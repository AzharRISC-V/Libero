`timescale 1 ns/100 ps
// Version: v12.2 12.700.0.21


module LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM(
       W_DATA,
       R_DATA,
       W_ADDR,
       R_ADDR,
       W_EN,
       R_EN,
       CLK,
       WBYTE_EN
    );
input  [79:0] W_DATA;
output [79:0] R_DATA;
input  [12:0] W_ADDR;
input  [12:0] R_ADDR;
input  W_EN;
input  R_EN;
input  CLK;
input  [7:0] WBYTE_EN;

    wire \R_DATA_TEMPR0[0] , \R_DATA_TEMPR1[0] , \R_DATA_TEMPR2[0] , 
        \R_DATA_TEMPR3[0] , \R_DATA_TEMPR4[0] , \R_DATA_TEMPR5[0] , 
        \R_DATA_TEMPR6[0] , \R_DATA_TEMPR7[0] , \R_DATA_TEMPR8[0] , 
        \R_DATA_TEMPR9[0] , \R_DATA_TEMPR10[0] , \R_DATA_TEMPR11[0] , 
        \R_DATA_TEMPR12[0] , \R_DATA_TEMPR13[0] , \R_DATA_TEMPR14[0] , 
        \R_DATA_TEMPR15[0] , \R_DATA_TEMPR0[1] , \R_DATA_TEMPR1[1] , 
        \R_DATA_TEMPR2[1] , \R_DATA_TEMPR3[1] , \R_DATA_TEMPR4[1] , 
        \R_DATA_TEMPR5[1] , \R_DATA_TEMPR6[1] , \R_DATA_TEMPR7[1] , 
        \R_DATA_TEMPR8[1] , \R_DATA_TEMPR9[1] , \R_DATA_TEMPR10[1] , 
        \R_DATA_TEMPR11[1] , \R_DATA_TEMPR12[1] , \R_DATA_TEMPR13[1] , 
        \R_DATA_TEMPR14[1] , \R_DATA_TEMPR15[1] , \R_DATA_TEMPR0[2] , 
        \R_DATA_TEMPR1[2] , \R_DATA_TEMPR2[2] , \R_DATA_TEMPR3[2] , 
        \R_DATA_TEMPR4[2] , \R_DATA_TEMPR5[2] , \R_DATA_TEMPR6[2] , 
        \R_DATA_TEMPR7[2] , \R_DATA_TEMPR8[2] , \R_DATA_TEMPR9[2] , 
        \R_DATA_TEMPR10[2] , \R_DATA_TEMPR11[2] , \R_DATA_TEMPR12[2] , 
        \R_DATA_TEMPR13[2] , \R_DATA_TEMPR14[2] , \R_DATA_TEMPR15[2] , 
        \R_DATA_TEMPR0[3] , \R_DATA_TEMPR1[3] , \R_DATA_TEMPR2[3] , 
        \R_DATA_TEMPR3[3] , \R_DATA_TEMPR4[3] , \R_DATA_TEMPR5[3] , 
        \R_DATA_TEMPR6[3] , \R_DATA_TEMPR7[3] , \R_DATA_TEMPR8[3] , 
        \R_DATA_TEMPR9[3] , \R_DATA_TEMPR10[3] , \R_DATA_TEMPR11[3] , 
        \R_DATA_TEMPR12[3] , \R_DATA_TEMPR13[3] , \R_DATA_TEMPR14[3] , 
        \R_DATA_TEMPR15[3] , \R_DATA_TEMPR0[4] , \R_DATA_TEMPR1[4] , 
        \R_DATA_TEMPR2[4] , \R_DATA_TEMPR3[4] , \R_DATA_TEMPR4[4] , 
        \R_DATA_TEMPR5[4] , \R_DATA_TEMPR6[4] , \R_DATA_TEMPR7[4] , 
        \R_DATA_TEMPR8[4] , \R_DATA_TEMPR9[4] , \R_DATA_TEMPR10[4] , 
        \R_DATA_TEMPR11[4] , \R_DATA_TEMPR12[4] , \R_DATA_TEMPR13[4] , 
        \R_DATA_TEMPR14[4] , \R_DATA_TEMPR15[4] , \R_DATA_TEMPR0[5] , 
        \R_DATA_TEMPR1[5] , \R_DATA_TEMPR2[5] , \R_DATA_TEMPR3[5] , 
        \R_DATA_TEMPR4[5] , \R_DATA_TEMPR5[5] , \R_DATA_TEMPR6[5] , 
        \R_DATA_TEMPR7[5] , \R_DATA_TEMPR8[5] , \R_DATA_TEMPR9[5] , 
        \R_DATA_TEMPR10[5] , \R_DATA_TEMPR11[5] , \R_DATA_TEMPR12[5] , 
        \R_DATA_TEMPR13[5] , \R_DATA_TEMPR14[5] , \R_DATA_TEMPR15[5] , 
        \R_DATA_TEMPR0[6] , \R_DATA_TEMPR1[6] , \R_DATA_TEMPR2[6] , 
        \R_DATA_TEMPR3[6] , \R_DATA_TEMPR4[6] , \R_DATA_TEMPR5[6] , 
        \R_DATA_TEMPR6[6] , \R_DATA_TEMPR7[6] , \R_DATA_TEMPR8[6] , 
        \R_DATA_TEMPR9[6] , \R_DATA_TEMPR10[6] , \R_DATA_TEMPR11[6] , 
        \R_DATA_TEMPR12[6] , \R_DATA_TEMPR13[6] , \R_DATA_TEMPR14[6] , 
        \R_DATA_TEMPR15[6] , \R_DATA_TEMPR0[7] , \R_DATA_TEMPR1[7] , 
        \R_DATA_TEMPR2[7] , \R_DATA_TEMPR3[7] , \R_DATA_TEMPR4[7] , 
        \R_DATA_TEMPR5[7] , \R_DATA_TEMPR6[7] , \R_DATA_TEMPR7[7] , 
        \R_DATA_TEMPR8[7] , \R_DATA_TEMPR9[7] , \R_DATA_TEMPR10[7] , 
        \R_DATA_TEMPR11[7] , \R_DATA_TEMPR12[7] , \R_DATA_TEMPR13[7] , 
        \R_DATA_TEMPR14[7] , \R_DATA_TEMPR15[7] , \R_DATA_TEMPR0[8] , 
        \R_DATA_TEMPR1[8] , \R_DATA_TEMPR2[8] , \R_DATA_TEMPR3[8] , 
        \R_DATA_TEMPR4[8] , \R_DATA_TEMPR5[8] , \R_DATA_TEMPR6[8] , 
        \R_DATA_TEMPR7[8] , \R_DATA_TEMPR8[8] , \R_DATA_TEMPR9[8] , 
        \R_DATA_TEMPR10[8] , \R_DATA_TEMPR11[8] , \R_DATA_TEMPR12[8] , 
        \R_DATA_TEMPR13[8] , \R_DATA_TEMPR14[8] , \R_DATA_TEMPR15[8] , 
        \R_DATA_TEMPR0[9] , \R_DATA_TEMPR1[9] , \R_DATA_TEMPR2[9] , 
        \R_DATA_TEMPR3[9] , \R_DATA_TEMPR4[9] , \R_DATA_TEMPR5[9] , 
        \R_DATA_TEMPR6[9] , \R_DATA_TEMPR7[9] , \R_DATA_TEMPR8[9] , 
        \R_DATA_TEMPR9[9] , \R_DATA_TEMPR10[9] , \R_DATA_TEMPR11[9] , 
        \R_DATA_TEMPR12[9] , \R_DATA_TEMPR13[9] , \R_DATA_TEMPR14[9] , 
        \R_DATA_TEMPR15[9] , \R_DATA_TEMPR0[10] , \R_DATA_TEMPR1[10] , 
        \R_DATA_TEMPR2[10] , \R_DATA_TEMPR3[10] , \R_DATA_TEMPR4[10] , 
        \R_DATA_TEMPR5[10] , \R_DATA_TEMPR6[10] , \R_DATA_TEMPR7[10] , 
        \R_DATA_TEMPR8[10] , \R_DATA_TEMPR9[10] , \R_DATA_TEMPR10[10] , 
        \R_DATA_TEMPR11[10] , \R_DATA_TEMPR12[10] , 
        \R_DATA_TEMPR13[10] , \R_DATA_TEMPR14[10] , 
        \R_DATA_TEMPR15[10] , \R_DATA_TEMPR0[11] , \R_DATA_TEMPR1[11] , 
        \R_DATA_TEMPR2[11] , \R_DATA_TEMPR3[11] , \R_DATA_TEMPR4[11] , 
        \R_DATA_TEMPR5[11] , \R_DATA_TEMPR6[11] , \R_DATA_TEMPR7[11] , 
        \R_DATA_TEMPR8[11] , \R_DATA_TEMPR9[11] , \R_DATA_TEMPR10[11] , 
        \R_DATA_TEMPR11[11] , \R_DATA_TEMPR12[11] , 
        \R_DATA_TEMPR13[11] , \R_DATA_TEMPR14[11] , 
        \R_DATA_TEMPR15[11] , \R_DATA_TEMPR0[12] , \R_DATA_TEMPR1[12] , 
        \R_DATA_TEMPR2[12] , \R_DATA_TEMPR3[12] , \R_DATA_TEMPR4[12] , 
        \R_DATA_TEMPR5[12] , \R_DATA_TEMPR6[12] , \R_DATA_TEMPR7[12] , 
        \R_DATA_TEMPR8[12] , \R_DATA_TEMPR9[12] , \R_DATA_TEMPR10[12] , 
        \R_DATA_TEMPR11[12] , \R_DATA_TEMPR12[12] , 
        \R_DATA_TEMPR13[12] , \R_DATA_TEMPR14[12] , 
        \R_DATA_TEMPR15[12] , \R_DATA_TEMPR0[13] , \R_DATA_TEMPR1[13] , 
        \R_DATA_TEMPR2[13] , \R_DATA_TEMPR3[13] , \R_DATA_TEMPR4[13] , 
        \R_DATA_TEMPR5[13] , \R_DATA_TEMPR6[13] , \R_DATA_TEMPR7[13] , 
        \R_DATA_TEMPR8[13] , \R_DATA_TEMPR9[13] , \R_DATA_TEMPR10[13] , 
        \R_DATA_TEMPR11[13] , \R_DATA_TEMPR12[13] , 
        \R_DATA_TEMPR13[13] , \R_DATA_TEMPR14[13] , 
        \R_DATA_TEMPR15[13] , \R_DATA_TEMPR0[14] , \R_DATA_TEMPR1[14] , 
        \R_DATA_TEMPR2[14] , \R_DATA_TEMPR3[14] , \R_DATA_TEMPR4[14] , 
        \R_DATA_TEMPR5[14] , \R_DATA_TEMPR6[14] , \R_DATA_TEMPR7[14] , 
        \R_DATA_TEMPR8[14] , \R_DATA_TEMPR9[14] , \R_DATA_TEMPR10[14] , 
        \R_DATA_TEMPR11[14] , \R_DATA_TEMPR12[14] , 
        \R_DATA_TEMPR13[14] , \R_DATA_TEMPR14[14] , 
        \R_DATA_TEMPR15[14] , \R_DATA_TEMPR0[15] , \R_DATA_TEMPR1[15] , 
        \R_DATA_TEMPR2[15] , \R_DATA_TEMPR3[15] , \R_DATA_TEMPR4[15] , 
        \R_DATA_TEMPR5[15] , \R_DATA_TEMPR6[15] , \R_DATA_TEMPR7[15] , 
        \R_DATA_TEMPR8[15] , \R_DATA_TEMPR9[15] , \R_DATA_TEMPR10[15] , 
        \R_DATA_TEMPR11[15] , \R_DATA_TEMPR12[15] , 
        \R_DATA_TEMPR13[15] , \R_DATA_TEMPR14[15] , 
        \R_DATA_TEMPR15[15] , \R_DATA_TEMPR0[16] , \R_DATA_TEMPR1[16] , 
        \R_DATA_TEMPR2[16] , \R_DATA_TEMPR3[16] , \R_DATA_TEMPR4[16] , 
        \R_DATA_TEMPR5[16] , \R_DATA_TEMPR6[16] , \R_DATA_TEMPR7[16] , 
        \R_DATA_TEMPR8[16] , \R_DATA_TEMPR9[16] , \R_DATA_TEMPR10[16] , 
        \R_DATA_TEMPR11[16] , \R_DATA_TEMPR12[16] , 
        \R_DATA_TEMPR13[16] , \R_DATA_TEMPR14[16] , 
        \R_DATA_TEMPR15[16] , \R_DATA_TEMPR0[17] , \R_DATA_TEMPR1[17] , 
        \R_DATA_TEMPR2[17] , \R_DATA_TEMPR3[17] , \R_DATA_TEMPR4[17] , 
        \R_DATA_TEMPR5[17] , \R_DATA_TEMPR6[17] , \R_DATA_TEMPR7[17] , 
        \R_DATA_TEMPR8[17] , \R_DATA_TEMPR9[17] , \R_DATA_TEMPR10[17] , 
        \R_DATA_TEMPR11[17] , \R_DATA_TEMPR12[17] , 
        \R_DATA_TEMPR13[17] , \R_DATA_TEMPR14[17] , 
        \R_DATA_TEMPR15[17] , \R_DATA_TEMPR0[18] , \R_DATA_TEMPR1[18] , 
        \R_DATA_TEMPR2[18] , \R_DATA_TEMPR3[18] , \R_DATA_TEMPR4[18] , 
        \R_DATA_TEMPR5[18] , \R_DATA_TEMPR6[18] , \R_DATA_TEMPR7[18] , 
        \R_DATA_TEMPR8[18] , \R_DATA_TEMPR9[18] , \R_DATA_TEMPR10[18] , 
        \R_DATA_TEMPR11[18] , \R_DATA_TEMPR12[18] , 
        \R_DATA_TEMPR13[18] , \R_DATA_TEMPR14[18] , 
        \R_DATA_TEMPR15[18] , \R_DATA_TEMPR0[19] , \R_DATA_TEMPR1[19] , 
        \R_DATA_TEMPR2[19] , \R_DATA_TEMPR3[19] , \R_DATA_TEMPR4[19] , 
        \R_DATA_TEMPR5[19] , \R_DATA_TEMPR6[19] , \R_DATA_TEMPR7[19] , 
        \R_DATA_TEMPR8[19] , \R_DATA_TEMPR9[19] , \R_DATA_TEMPR10[19] , 
        \R_DATA_TEMPR11[19] , \R_DATA_TEMPR12[19] , 
        \R_DATA_TEMPR13[19] , \R_DATA_TEMPR14[19] , 
        \R_DATA_TEMPR15[19] , \R_DATA_TEMPR0[20] , \R_DATA_TEMPR1[20] , 
        \R_DATA_TEMPR2[20] , \R_DATA_TEMPR3[20] , \R_DATA_TEMPR4[20] , 
        \R_DATA_TEMPR5[20] , \R_DATA_TEMPR6[20] , \R_DATA_TEMPR7[20] , 
        \R_DATA_TEMPR8[20] , \R_DATA_TEMPR9[20] , \R_DATA_TEMPR10[20] , 
        \R_DATA_TEMPR11[20] , \R_DATA_TEMPR12[20] , 
        \R_DATA_TEMPR13[20] , \R_DATA_TEMPR14[20] , 
        \R_DATA_TEMPR15[20] , \R_DATA_TEMPR0[21] , \R_DATA_TEMPR1[21] , 
        \R_DATA_TEMPR2[21] , \R_DATA_TEMPR3[21] , \R_DATA_TEMPR4[21] , 
        \R_DATA_TEMPR5[21] , \R_DATA_TEMPR6[21] , \R_DATA_TEMPR7[21] , 
        \R_DATA_TEMPR8[21] , \R_DATA_TEMPR9[21] , \R_DATA_TEMPR10[21] , 
        \R_DATA_TEMPR11[21] , \R_DATA_TEMPR12[21] , 
        \R_DATA_TEMPR13[21] , \R_DATA_TEMPR14[21] , 
        \R_DATA_TEMPR15[21] , \R_DATA_TEMPR0[22] , \R_DATA_TEMPR1[22] , 
        \R_DATA_TEMPR2[22] , \R_DATA_TEMPR3[22] , \R_DATA_TEMPR4[22] , 
        \R_DATA_TEMPR5[22] , \R_DATA_TEMPR6[22] , \R_DATA_TEMPR7[22] , 
        \R_DATA_TEMPR8[22] , \R_DATA_TEMPR9[22] , \R_DATA_TEMPR10[22] , 
        \R_DATA_TEMPR11[22] , \R_DATA_TEMPR12[22] , 
        \R_DATA_TEMPR13[22] , \R_DATA_TEMPR14[22] , 
        \R_DATA_TEMPR15[22] , \R_DATA_TEMPR0[23] , \R_DATA_TEMPR1[23] , 
        \R_DATA_TEMPR2[23] , \R_DATA_TEMPR3[23] , \R_DATA_TEMPR4[23] , 
        \R_DATA_TEMPR5[23] , \R_DATA_TEMPR6[23] , \R_DATA_TEMPR7[23] , 
        \R_DATA_TEMPR8[23] , \R_DATA_TEMPR9[23] , \R_DATA_TEMPR10[23] , 
        \R_DATA_TEMPR11[23] , \R_DATA_TEMPR12[23] , 
        \R_DATA_TEMPR13[23] , \R_DATA_TEMPR14[23] , 
        \R_DATA_TEMPR15[23] , \R_DATA_TEMPR0[24] , \R_DATA_TEMPR1[24] , 
        \R_DATA_TEMPR2[24] , \R_DATA_TEMPR3[24] , \R_DATA_TEMPR4[24] , 
        \R_DATA_TEMPR5[24] , \R_DATA_TEMPR6[24] , \R_DATA_TEMPR7[24] , 
        \R_DATA_TEMPR8[24] , \R_DATA_TEMPR9[24] , \R_DATA_TEMPR10[24] , 
        \R_DATA_TEMPR11[24] , \R_DATA_TEMPR12[24] , 
        \R_DATA_TEMPR13[24] , \R_DATA_TEMPR14[24] , 
        \R_DATA_TEMPR15[24] , \R_DATA_TEMPR0[25] , \R_DATA_TEMPR1[25] , 
        \R_DATA_TEMPR2[25] , \R_DATA_TEMPR3[25] , \R_DATA_TEMPR4[25] , 
        \R_DATA_TEMPR5[25] , \R_DATA_TEMPR6[25] , \R_DATA_TEMPR7[25] , 
        \R_DATA_TEMPR8[25] , \R_DATA_TEMPR9[25] , \R_DATA_TEMPR10[25] , 
        \R_DATA_TEMPR11[25] , \R_DATA_TEMPR12[25] , 
        \R_DATA_TEMPR13[25] , \R_DATA_TEMPR14[25] , 
        \R_DATA_TEMPR15[25] , \R_DATA_TEMPR0[26] , \R_DATA_TEMPR1[26] , 
        \R_DATA_TEMPR2[26] , \R_DATA_TEMPR3[26] , \R_DATA_TEMPR4[26] , 
        \R_DATA_TEMPR5[26] , \R_DATA_TEMPR6[26] , \R_DATA_TEMPR7[26] , 
        \R_DATA_TEMPR8[26] , \R_DATA_TEMPR9[26] , \R_DATA_TEMPR10[26] , 
        \R_DATA_TEMPR11[26] , \R_DATA_TEMPR12[26] , 
        \R_DATA_TEMPR13[26] , \R_DATA_TEMPR14[26] , 
        \R_DATA_TEMPR15[26] , \R_DATA_TEMPR0[27] , \R_DATA_TEMPR1[27] , 
        \R_DATA_TEMPR2[27] , \R_DATA_TEMPR3[27] , \R_DATA_TEMPR4[27] , 
        \R_DATA_TEMPR5[27] , \R_DATA_TEMPR6[27] , \R_DATA_TEMPR7[27] , 
        \R_DATA_TEMPR8[27] , \R_DATA_TEMPR9[27] , \R_DATA_TEMPR10[27] , 
        \R_DATA_TEMPR11[27] , \R_DATA_TEMPR12[27] , 
        \R_DATA_TEMPR13[27] , \R_DATA_TEMPR14[27] , 
        \R_DATA_TEMPR15[27] , \R_DATA_TEMPR0[28] , \R_DATA_TEMPR1[28] , 
        \R_DATA_TEMPR2[28] , \R_DATA_TEMPR3[28] , \R_DATA_TEMPR4[28] , 
        \R_DATA_TEMPR5[28] , \R_DATA_TEMPR6[28] , \R_DATA_TEMPR7[28] , 
        \R_DATA_TEMPR8[28] , \R_DATA_TEMPR9[28] , \R_DATA_TEMPR10[28] , 
        \R_DATA_TEMPR11[28] , \R_DATA_TEMPR12[28] , 
        \R_DATA_TEMPR13[28] , \R_DATA_TEMPR14[28] , 
        \R_DATA_TEMPR15[28] , \R_DATA_TEMPR0[29] , \R_DATA_TEMPR1[29] , 
        \R_DATA_TEMPR2[29] , \R_DATA_TEMPR3[29] , \R_DATA_TEMPR4[29] , 
        \R_DATA_TEMPR5[29] , \R_DATA_TEMPR6[29] , \R_DATA_TEMPR7[29] , 
        \R_DATA_TEMPR8[29] , \R_DATA_TEMPR9[29] , \R_DATA_TEMPR10[29] , 
        \R_DATA_TEMPR11[29] , \R_DATA_TEMPR12[29] , 
        \R_DATA_TEMPR13[29] , \R_DATA_TEMPR14[29] , 
        \R_DATA_TEMPR15[29] , \R_DATA_TEMPR0[30] , \R_DATA_TEMPR1[30] , 
        \R_DATA_TEMPR2[30] , \R_DATA_TEMPR3[30] , \R_DATA_TEMPR4[30] , 
        \R_DATA_TEMPR5[30] , \R_DATA_TEMPR6[30] , \R_DATA_TEMPR7[30] , 
        \R_DATA_TEMPR8[30] , \R_DATA_TEMPR9[30] , \R_DATA_TEMPR10[30] , 
        \R_DATA_TEMPR11[30] , \R_DATA_TEMPR12[30] , 
        \R_DATA_TEMPR13[30] , \R_DATA_TEMPR14[30] , 
        \R_DATA_TEMPR15[30] , \R_DATA_TEMPR0[31] , \R_DATA_TEMPR1[31] , 
        \R_DATA_TEMPR2[31] , \R_DATA_TEMPR3[31] , \R_DATA_TEMPR4[31] , 
        \R_DATA_TEMPR5[31] , \R_DATA_TEMPR6[31] , \R_DATA_TEMPR7[31] , 
        \R_DATA_TEMPR8[31] , \R_DATA_TEMPR9[31] , \R_DATA_TEMPR10[31] , 
        \R_DATA_TEMPR11[31] , \R_DATA_TEMPR12[31] , 
        \R_DATA_TEMPR13[31] , \R_DATA_TEMPR14[31] , 
        \R_DATA_TEMPR15[31] , \R_DATA_TEMPR0[32] , \R_DATA_TEMPR1[32] , 
        \R_DATA_TEMPR2[32] , \R_DATA_TEMPR3[32] , \R_DATA_TEMPR4[32] , 
        \R_DATA_TEMPR5[32] , \R_DATA_TEMPR6[32] , \R_DATA_TEMPR7[32] , 
        \R_DATA_TEMPR8[32] , \R_DATA_TEMPR9[32] , \R_DATA_TEMPR10[32] , 
        \R_DATA_TEMPR11[32] , \R_DATA_TEMPR12[32] , 
        \R_DATA_TEMPR13[32] , \R_DATA_TEMPR14[32] , 
        \R_DATA_TEMPR15[32] , \R_DATA_TEMPR0[33] , \R_DATA_TEMPR1[33] , 
        \R_DATA_TEMPR2[33] , \R_DATA_TEMPR3[33] , \R_DATA_TEMPR4[33] , 
        \R_DATA_TEMPR5[33] , \R_DATA_TEMPR6[33] , \R_DATA_TEMPR7[33] , 
        \R_DATA_TEMPR8[33] , \R_DATA_TEMPR9[33] , \R_DATA_TEMPR10[33] , 
        \R_DATA_TEMPR11[33] , \R_DATA_TEMPR12[33] , 
        \R_DATA_TEMPR13[33] , \R_DATA_TEMPR14[33] , 
        \R_DATA_TEMPR15[33] , \R_DATA_TEMPR0[34] , \R_DATA_TEMPR1[34] , 
        \R_DATA_TEMPR2[34] , \R_DATA_TEMPR3[34] , \R_DATA_TEMPR4[34] , 
        \R_DATA_TEMPR5[34] , \R_DATA_TEMPR6[34] , \R_DATA_TEMPR7[34] , 
        \R_DATA_TEMPR8[34] , \R_DATA_TEMPR9[34] , \R_DATA_TEMPR10[34] , 
        \R_DATA_TEMPR11[34] , \R_DATA_TEMPR12[34] , 
        \R_DATA_TEMPR13[34] , \R_DATA_TEMPR14[34] , 
        \R_DATA_TEMPR15[34] , \R_DATA_TEMPR0[35] , \R_DATA_TEMPR1[35] , 
        \R_DATA_TEMPR2[35] , \R_DATA_TEMPR3[35] , \R_DATA_TEMPR4[35] , 
        \R_DATA_TEMPR5[35] , \R_DATA_TEMPR6[35] , \R_DATA_TEMPR7[35] , 
        \R_DATA_TEMPR8[35] , \R_DATA_TEMPR9[35] , \R_DATA_TEMPR10[35] , 
        \R_DATA_TEMPR11[35] , \R_DATA_TEMPR12[35] , 
        \R_DATA_TEMPR13[35] , \R_DATA_TEMPR14[35] , 
        \R_DATA_TEMPR15[35] , \R_DATA_TEMPR0[36] , \R_DATA_TEMPR1[36] , 
        \R_DATA_TEMPR2[36] , \R_DATA_TEMPR3[36] , \R_DATA_TEMPR4[36] , 
        \R_DATA_TEMPR5[36] , \R_DATA_TEMPR6[36] , \R_DATA_TEMPR7[36] , 
        \R_DATA_TEMPR8[36] , \R_DATA_TEMPR9[36] , \R_DATA_TEMPR10[36] , 
        \R_DATA_TEMPR11[36] , \R_DATA_TEMPR12[36] , 
        \R_DATA_TEMPR13[36] , \R_DATA_TEMPR14[36] , 
        \R_DATA_TEMPR15[36] , \R_DATA_TEMPR0[37] , \R_DATA_TEMPR1[37] , 
        \R_DATA_TEMPR2[37] , \R_DATA_TEMPR3[37] , \R_DATA_TEMPR4[37] , 
        \R_DATA_TEMPR5[37] , \R_DATA_TEMPR6[37] , \R_DATA_TEMPR7[37] , 
        \R_DATA_TEMPR8[37] , \R_DATA_TEMPR9[37] , \R_DATA_TEMPR10[37] , 
        \R_DATA_TEMPR11[37] , \R_DATA_TEMPR12[37] , 
        \R_DATA_TEMPR13[37] , \R_DATA_TEMPR14[37] , 
        \R_DATA_TEMPR15[37] , \R_DATA_TEMPR0[38] , \R_DATA_TEMPR1[38] , 
        \R_DATA_TEMPR2[38] , \R_DATA_TEMPR3[38] , \R_DATA_TEMPR4[38] , 
        \R_DATA_TEMPR5[38] , \R_DATA_TEMPR6[38] , \R_DATA_TEMPR7[38] , 
        \R_DATA_TEMPR8[38] , \R_DATA_TEMPR9[38] , \R_DATA_TEMPR10[38] , 
        \R_DATA_TEMPR11[38] , \R_DATA_TEMPR12[38] , 
        \R_DATA_TEMPR13[38] , \R_DATA_TEMPR14[38] , 
        \R_DATA_TEMPR15[38] , \R_DATA_TEMPR0[39] , \R_DATA_TEMPR1[39] , 
        \R_DATA_TEMPR2[39] , \R_DATA_TEMPR3[39] , \R_DATA_TEMPR4[39] , 
        \R_DATA_TEMPR5[39] , \R_DATA_TEMPR6[39] , \R_DATA_TEMPR7[39] , 
        \R_DATA_TEMPR8[39] , \R_DATA_TEMPR9[39] , \R_DATA_TEMPR10[39] , 
        \R_DATA_TEMPR11[39] , \R_DATA_TEMPR12[39] , 
        \R_DATA_TEMPR13[39] , \R_DATA_TEMPR14[39] , 
        \R_DATA_TEMPR15[39] , \R_DATA_TEMPR0[40] , \R_DATA_TEMPR1[40] , 
        \R_DATA_TEMPR2[40] , \R_DATA_TEMPR3[40] , \R_DATA_TEMPR4[40] , 
        \R_DATA_TEMPR5[40] , \R_DATA_TEMPR6[40] , \R_DATA_TEMPR7[40] , 
        \R_DATA_TEMPR8[40] , \R_DATA_TEMPR9[40] , \R_DATA_TEMPR10[40] , 
        \R_DATA_TEMPR11[40] , \R_DATA_TEMPR12[40] , 
        \R_DATA_TEMPR13[40] , \R_DATA_TEMPR14[40] , 
        \R_DATA_TEMPR15[40] , \R_DATA_TEMPR0[41] , \R_DATA_TEMPR1[41] , 
        \R_DATA_TEMPR2[41] , \R_DATA_TEMPR3[41] , \R_DATA_TEMPR4[41] , 
        \R_DATA_TEMPR5[41] , \R_DATA_TEMPR6[41] , \R_DATA_TEMPR7[41] , 
        \R_DATA_TEMPR8[41] , \R_DATA_TEMPR9[41] , \R_DATA_TEMPR10[41] , 
        \R_DATA_TEMPR11[41] , \R_DATA_TEMPR12[41] , 
        \R_DATA_TEMPR13[41] , \R_DATA_TEMPR14[41] , 
        \R_DATA_TEMPR15[41] , \R_DATA_TEMPR0[42] , \R_DATA_TEMPR1[42] , 
        \R_DATA_TEMPR2[42] , \R_DATA_TEMPR3[42] , \R_DATA_TEMPR4[42] , 
        \R_DATA_TEMPR5[42] , \R_DATA_TEMPR6[42] , \R_DATA_TEMPR7[42] , 
        \R_DATA_TEMPR8[42] , \R_DATA_TEMPR9[42] , \R_DATA_TEMPR10[42] , 
        \R_DATA_TEMPR11[42] , \R_DATA_TEMPR12[42] , 
        \R_DATA_TEMPR13[42] , \R_DATA_TEMPR14[42] , 
        \R_DATA_TEMPR15[42] , \R_DATA_TEMPR0[43] , \R_DATA_TEMPR1[43] , 
        \R_DATA_TEMPR2[43] , \R_DATA_TEMPR3[43] , \R_DATA_TEMPR4[43] , 
        \R_DATA_TEMPR5[43] , \R_DATA_TEMPR6[43] , \R_DATA_TEMPR7[43] , 
        \R_DATA_TEMPR8[43] , \R_DATA_TEMPR9[43] , \R_DATA_TEMPR10[43] , 
        \R_DATA_TEMPR11[43] , \R_DATA_TEMPR12[43] , 
        \R_DATA_TEMPR13[43] , \R_DATA_TEMPR14[43] , 
        \R_DATA_TEMPR15[43] , \R_DATA_TEMPR0[44] , \R_DATA_TEMPR1[44] , 
        \R_DATA_TEMPR2[44] , \R_DATA_TEMPR3[44] , \R_DATA_TEMPR4[44] , 
        \R_DATA_TEMPR5[44] , \R_DATA_TEMPR6[44] , \R_DATA_TEMPR7[44] , 
        \R_DATA_TEMPR8[44] , \R_DATA_TEMPR9[44] , \R_DATA_TEMPR10[44] , 
        \R_DATA_TEMPR11[44] , \R_DATA_TEMPR12[44] , 
        \R_DATA_TEMPR13[44] , \R_DATA_TEMPR14[44] , 
        \R_DATA_TEMPR15[44] , \R_DATA_TEMPR0[45] , \R_DATA_TEMPR1[45] , 
        \R_DATA_TEMPR2[45] , \R_DATA_TEMPR3[45] , \R_DATA_TEMPR4[45] , 
        \R_DATA_TEMPR5[45] , \R_DATA_TEMPR6[45] , \R_DATA_TEMPR7[45] , 
        \R_DATA_TEMPR8[45] , \R_DATA_TEMPR9[45] , \R_DATA_TEMPR10[45] , 
        \R_DATA_TEMPR11[45] , \R_DATA_TEMPR12[45] , 
        \R_DATA_TEMPR13[45] , \R_DATA_TEMPR14[45] , 
        \R_DATA_TEMPR15[45] , \R_DATA_TEMPR0[46] , \R_DATA_TEMPR1[46] , 
        \R_DATA_TEMPR2[46] , \R_DATA_TEMPR3[46] , \R_DATA_TEMPR4[46] , 
        \R_DATA_TEMPR5[46] , \R_DATA_TEMPR6[46] , \R_DATA_TEMPR7[46] , 
        \R_DATA_TEMPR8[46] , \R_DATA_TEMPR9[46] , \R_DATA_TEMPR10[46] , 
        \R_DATA_TEMPR11[46] , \R_DATA_TEMPR12[46] , 
        \R_DATA_TEMPR13[46] , \R_DATA_TEMPR14[46] , 
        \R_DATA_TEMPR15[46] , \R_DATA_TEMPR0[47] , \R_DATA_TEMPR1[47] , 
        \R_DATA_TEMPR2[47] , \R_DATA_TEMPR3[47] , \R_DATA_TEMPR4[47] , 
        \R_DATA_TEMPR5[47] , \R_DATA_TEMPR6[47] , \R_DATA_TEMPR7[47] , 
        \R_DATA_TEMPR8[47] , \R_DATA_TEMPR9[47] , \R_DATA_TEMPR10[47] , 
        \R_DATA_TEMPR11[47] , \R_DATA_TEMPR12[47] , 
        \R_DATA_TEMPR13[47] , \R_DATA_TEMPR14[47] , 
        \R_DATA_TEMPR15[47] , \R_DATA_TEMPR0[48] , \R_DATA_TEMPR1[48] , 
        \R_DATA_TEMPR2[48] , \R_DATA_TEMPR3[48] , \R_DATA_TEMPR4[48] , 
        \R_DATA_TEMPR5[48] , \R_DATA_TEMPR6[48] , \R_DATA_TEMPR7[48] , 
        \R_DATA_TEMPR8[48] , \R_DATA_TEMPR9[48] , \R_DATA_TEMPR10[48] , 
        \R_DATA_TEMPR11[48] , \R_DATA_TEMPR12[48] , 
        \R_DATA_TEMPR13[48] , \R_DATA_TEMPR14[48] , 
        \R_DATA_TEMPR15[48] , \R_DATA_TEMPR0[49] , \R_DATA_TEMPR1[49] , 
        \R_DATA_TEMPR2[49] , \R_DATA_TEMPR3[49] , \R_DATA_TEMPR4[49] , 
        \R_DATA_TEMPR5[49] , \R_DATA_TEMPR6[49] , \R_DATA_TEMPR7[49] , 
        \R_DATA_TEMPR8[49] , \R_DATA_TEMPR9[49] , \R_DATA_TEMPR10[49] , 
        \R_DATA_TEMPR11[49] , \R_DATA_TEMPR12[49] , 
        \R_DATA_TEMPR13[49] , \R_DATA_TEMPR14[49] , 
        \R_DATA_TEMPR15[49] , \R_DATA_TEMPR0[50] , \R_DATA_TEMPR1[50] , 
        \R_DATA_TEMPR2[50] , \R_DATA_TEMPR3[50] , \R_DATA_TEMPR4[50] , 
        \R_DATA_TEMPR5[50] , \R_DATA_TEMPR6[50] , \R_DATA_TEMPR7[50] , 
        \R_DATA_TEMPR8[50] , \R_DATA_TEMPR9[50] , \R_DATA_TEMPR10[50] , 
        \R_DATA_TEMPR11[50] , \R_DATA_TEMPR12[50] , 
        \R_DATA_TEMPR13[50] , \R_DATA_TEMPR14[50] , 
        \R_DATA_TEMPR15[50] , \R_DATA_TEMPR0[51] , \R_DATA_TEMPR1[51] , 
        \R_DATA_TEMPR2[51] , \R_DATA_TEMPR3[51] , \R_DATA_TEMPR4[51] , 
        \R_DATA_TEMPR5[51] , \R_DATA_TEMPR6[51] , \R_DATA_TEMPR7[51] , 
        \R_DATA_TEMPR8[51] , \R_DATA_TEMPR9[51] , \R_DATA_TEMPR10[51] , 
        \R_DATA_TEMPR11[51] , \R_DATA_TEMPR12[51] , 
        \R_DATA_TEMPR13[51] , \R_DATA_TEMPR14[51] , 
        \R_DATA_TEMPR15[51] , \R_DATA_TEMPR0[52] , \R_DATA_TEMPR1[52] , 
        \R_DATA_TEMPR2[52] , \R_DATA_TEMPR3[52] , \R_DATA_TEMPR4[52] , 
        \R_DATA_TEMPR5[52] , \R_DATA_TEMPR6[52] , \R_DATA_TEMPR7[52] , 
        \R_DATA_TEMPR8[52] , \R_DATA_TEMPR9[52] , \R_DATA_TEMPR10[52] , 
        \R_DATA_TEMPR11[52] , \R_DATA_TEMPR12[52] , 
        \R_DATA_TEMPR13[52] , \R_DATA_TEMPR14[52] , 
        \R_DATA_TEMPR15[52] , \R_DATA_TEMPR0[53] , \R_DATA_TEMPR1[53] , 
        \R_DATA_TEMPR2[53] , \R_DATA_TEMPR3[53] , \R_DATA_TEMPR4[53] , 
        \R_DATA_TEMPR5[53] , \R_DATA_TEMPR6[53] , \R_DATA_TEMPR7[53] , 
        \R_DATA_TEMPR8[53] , \R_DATA_TEMPR9[53] , \R_DATA_TEMPR10[53] , 
        \R_DATA_TEMPR11[53] , \R_DATA_TEMPR12[53] , 
        \R_DATA_TEMPR13[53] , \R_DATA_TEMPR14[53] , 
        \R_DATA_TEMPR15[53] , \R_DATA_TEMPR0[54] , \R_DATA_TEMPR1[54] , 
        \R_DATA_TEMPR2[54] , \R_DATA_TEMPR3[54] , \R_DATA_TEMPR4[54] , 
        \R_DATA_TEMPR5[54] , \R_DATA_TEMPR6[54] , \R_DATA_TEMPR7[54] , 
        \R_DATA_TEMPR8[54] , \R_DATA_TEMPR9[54] , \R_DATA_TEMPR10[54] , 
        \R_DATA_TEMPR11[54] , \R_DATA_TEMPR12[54] , 
        \R_DATA_TEMPR13[54] , \R_DATA_TEMPR14[54] , 
        \R_DATA_TEMPR15[54] , \R_DATA_TEMPR0[55] , \R_DATA_TEMPR1[55] , 
        \R_DATA_TEMPR2[55] , \R_DATA_TEMPR3[55] , \R_DATA_TEMPR4[55] , 
        \R_DATA_TEMPR5[55] , \R_DATA_TEMPR6[55] , \R_DATA_TEMPR7[55] , 
        \R_DATA_TEMPR8[55] , \R_DATA_TEMPR9[55] , \R_DATA_TEMPR10[55] , 
        \R_DATA_TEMPR11[55] , \R_DATA_TEMPR12[55] , 
        \R_DATA_TEMPR13[55] , \R_DATA_TEMPR14[55] , 
        \R_DATA_TEMPR15[55] , \R_DATA_TEMPR0[56] , \R_DATA_TEMPR1[56] , 
        \R_DATA_TEMPR2[56] , \R_DATA_TEMPR3[56] , \R_DATA_TEMPR4[56] , 
        \R_DATA_TEMPR5[56] , \R_DATA_TEMPR6[56] , \R_DATA_TEMPR7[56] , 
        \R_DATA_TEMPR8[56] , \R_DATA_TEMPR9[56] , \R_DATA_TEMPR10[56] , 
        \R_DATA_TEMPR11[56] , \R_DATA_TEMPR12[56] , 
        \R_DATA_TEMPR13[56] , \R_DATA_TEMPR14[56] , 
        \R_DATA_TEMPR15[56] , \R_DATA_TEMPR0[57] , \R_DATA_TEMPR1[57] , 
        \R_DATA_TEMPR2[57] , \R_DATA_TEMPR3[57] , \R_DATA_TEMPR4[57] , 
        \R_DATA_TEMPR5[57] , \R_DATA_TEMPR6[57] , \R_DATA_TEMPR7[57] , 
        \R_DATA_TEMPR8[57] , \R_DATA_TEMPR9[57] , \R_DATA_TEMPR10[57] , 
        \R_DATA_TEMPR11[57] , \R_DATA_TEMPR12[57] , 
        \R_DATA_TEMPR13[57] , \R_DATA_TEMPR14[57] , 
        \R_DATA_TEMPR15[57] , \R_DATA_TEMPR0[58] , \R_DATA_TEMPR1[58] , 
        \R_DATA_TEMPR2[58] , \R_DATA_TEMPR3[58] , \R_DATA_TEMPR4[58] , 
        \R_DATA_TEMPR5[58] , \R_DATA_TEMPR6[58] , \R_DATA_TEMPR7[58] , 
        \R_DATA_TEMPR8[58] , \R_DATA_TEMPR9[58] , \R_DATA_TEMPR10[58] , 
        \R_DATA_TEMPR11[58] , \R_DATA_TEMPR12[58] , 
        \R_DATA_TEMPR13[58] , \R_DATA_TEMPR14[58] , 
        \R_DATA_TEMPR15[58] , \R_DATA_TEMPR0[59] , \R_DATA_TEMPR1[59] , 
        \R_DATA_TEMPR2[59] , \R_DATA_TEMPR3[59] , \R_DATA_TEMPR4[59] , 
        \R_DATA_TEMPR5[59] , \R_DATA_TEMPR6[59] , \R_DATA_TEMPR7[59] , 
        \R_DATA_TEMPR8[59] , \R_DATA_TEMPR9[59] , \R_DATA_TEMPR10[59] , 
        \R_DATA_TEMPR11[59] , \R_DATA_TEMPR12[59] , 
        \R_DATA_TEMPR13[59] , \R_DATA_TEMPR14[59] , 
        \R_DATA_TEMPR15[59] , \R_DATA_TEMPR0[60] , \R_DATA_TEMPR1[60] , 
        \R_DATA_TEMPR2[60] , \R_DATA_TEMPR3[60] , \R_DATA_TEMPR4[60] , 
        \R_DATA_TEMPR5[60] , \R_DATA_TEMPR6[60] , \R_DATA_TEMPR7[60] , 
        \R_DATA_TEMPR8[60] , \R_DATA_TEMPR9[60] , \R_DATA_TEMPR10[60] , 
        \R_DATA_TEMPR11[60] , \R_DATA_TEMPR12[60] , 
        \R_DATA_TEMPR13[60] , \R_DATA_TEMPR14[60] , 
        \R_DATA_TEMPR15[60] , \R_DATA_TEMPR0[61] , \R_DATA_TEMPR1[61] , 
        \R_DATA_TEMPR2[61] , \R_DATA_TEMPR3[61] , \R_DATA_TEMPR4[61] , 
        \R_DATA_TEMPR5[61] , \R_DATA_TEMPR6[61] , \R_DATA_TEMPR7[61] , 
        \R_DATA_TEMPR8[61] , \R_DATA_TEMPR9[61] , \R_DATA_TEMPR10[61] , 
        \R_DATA_TEMPR11[61] , \R_DATA_TEMPR12[61] , 
        \R_DATA_TEMPR13[61] , \R_DATA_TEMPR14[61] , 
        \R_DATA_TEMPR15[61] , \R_DATA_TEMPR0[62] , \R_DATA_TEMPR1[62] , 
        \R_DATA_TEMPR2[62] , \R_DATA_TEMPR3[62] , \R_DATA_TEMPR4[62] , 
        \R_DATA_TEMPR5[62] , \R_DATA_TEMPR6[62] , \R_DATA_TEMPR7[62] , 
        \R_DATA_TEMPR8[62] , \R_DATA_TEMPR9[62] , \R_DATA_TEMPR10[62] , 
        \R_DATA_TEMPR11[62] , \R_DATA_TEMPR12[62] , 
        \R_DATA_TEMPR13[62] , \R_DATA_TEMPR14[62] , 
        \R_DATA_TEMPR15[62] , \R_DATA_TEMPR0[63] , \R_DATA_TEMPR1[63] , 
        \R_DATA_TEMPR2[63] , \R_DATA_TEMPR3[63] , \R_DATA_TEMPR4[63] , 
        \R_DATA_TEMPR5[63] , \R_DATA_TEMPR6[63] , \R_DATA_TEMPR7[63] , 
        \R_DATA_TEMPR8[63] , \R_DATA_TEMPR9[63] , \R_DATA_TEMPR10[63] , 
        \R_DATA_TEMPR11[63] , \R_DATA_TEMPR12[63] , 
        \R_DATA_TEMPR13[63] , \R_DATA_TEMPR14[63] , 
        \R_DATA_TEMPR15[63] , \R_DATA_TEMPR0[64] , \R_DATA_TEMPR1[64] , 
        \R_DATA_TEMPR2[64] , \R_DATA_TEMPR3[64] , \R_DATA_TEMPR4[64] , 
        \R_DATA_TEMPR5[64] , \R_DATA_TEMPR6[64] , \R_DATA_TEMPR7[64] , 
        \R_DATA_TEMPR8[64] , \R_DATA_TEMPR9[64] , \R_DATA_TEMPR10[64] , 
        \R_DATA_TEMPR11[64] , \R_DATA_TEMPR12[64] , 
        \R_DATA_TEMPR13[64] , \R_DATA_TEMPR14[64] , 
        \R_DATA_TEMPR15[64] , \R_DATA_TEMPR0[65] , \R_DATA_TEMPR1[65] , 
        \R_DATA_TEMPR2[65] , \R_DATA_TEMPR3[65] , \R_DATA_TEMPR4[65] , 
        \R_DATA_TEMPR5[65] , \R_DATA_TEMPR6[65] , \R_DATA_TEMPR7[65] , 
        \R_DATA_TEMPR8[65] , \R_DATA_TEMPR9[65] , \R_DATA_TEMPR10[65] , 
        \R_DATA_TEMPR11[65] , \R_DATA_TEMPR12[65] , 
        \R_DATA_TEMPR13[65] , \R_DATA_TEMPR14[65] , 
        \R_DATA_TEMPR15[65] , \R_DATA_TEMPR0[66] , \R_DATA_TEMPR1[66] , 
        \R_DATA_TEMPR2[66] , \R_DATA_TEMPR3[66] , \R_DATA_TEMPR4[66] , 
        \R_DATA_TEMPR5[66] , \R_DATA_TEMPR6[66] , \R_DATA_TEMPR7[66] , 
        \R_DATA_TEMPR8[66] , \R_DATA_TEMPR9[66] , \R_DATA_TEMPR10[66] , 
        \R_DATA_TEMPR11[66] , \R_DATA_TEMPR12[66] , 
        \R_DATA_TEMPR13[66] , \R_DATA_TEMPR14[66] , 
        \R_DATA_TEMPR15[66] , \R_DATA_TEMPR0[67] , \R_DATA_TEMPR1[67] , 
        \R_DATA_TEMPR2[67] , \R_DATA_TEMPR3[67] , \R_DATA_TEMPR4[67] , 
        \R_DATA_TEMPR5[67] , \R_DATA_TEMPR6[67] , \R_DATA_TEMPR7[67] , 
        \R_DATA_TEMPR8[67] , \R_DATA_TEMPR9[67] , \R_DATA_TEMPR10[67] , 
        \R_DATA_TEMPR11[67] , \R_DATA_TEMPR12[67] , 
        \R_DATA_TEMPR13[67] , \R_DATA_TEMPR14[67] , 
        \R_DATA_TEMPR15[67] , \R_DATA_TEMPR0[68] , \R_DATA_TEMPR1[68] , 
        \R_DATA_TEMPR2[68] , \R_DATA_TEMPR3[68] , \R_DATA_TEMPR4[68] , 
        \R_DATA_TEMPR5[68] , \R_DATA_TEMPR6[68] , \R_DATA_TEMPR7[68] , 
        \R_DATA_TEMPR8[68] , \R_DATA_TEMPR9[68] , \R_DATA_TEMPR10[68] , 
        \R_DATA_TEMPR11[68] , \R_DATA_TEMPR12[68] , 
        \R_DATA_TEMPR13[68] , \R_DATA_TEMPR14[68] , 
        \R_DATA_TEMPR15[68] , \R_DATA_TEMPR0[69] , \R_DATA_TEMPR1[69] , 
        \R_DATA_TEMPR2[69] , \R_DATA_TEMPR3[69] , \R_DATA_TEMPR4[69] , 
        \R_DATA_TEMPR5[69] , \R_DATA_TEMPR6[69] , \R_DATA_TEMPR7[69] , 
        \R_DATA_TEMPR8[69] , \R_DATA_TEMPR9[69] , \R_DATA_TEMPR10[69] , 
        \R_DATA_TEMPR11[69] , \R_DATA_TEMPR12[69] , 
        \R_DATA_TEMPR13[69] , \R_DATA_TEMPR14[69] , 
        \R_DATA_TEMPR15[69] , \R_DATA_TEMPR0[70] , \R_DATA_TEMPR1[70] , 
        \R_DATA_TEMPR2[70] , \R_DATA_TEMPR3[70] , \R_DATA_TEMPR4[70] , 
        \R_DATA_TEMPR5[70] , \R_DATA_TEMPR6[70] , \R_DATA_TEMPR7[70] , 
        \R_DATA_TEMPR8[70] , \R_DATA_TEMPR9[70] , \R_DATA_TEMPR10[70] , 
        \R_DATA_TEMPR11[70] , \R_DATA_TEMPR12[70] , 
        \R_DATA_TEMPR13[70] , \R_DATA_TEMPR14[70] , 
        \R_DATA_TEMPR15[70] , \R_DATA_TEMPR0[71] , \R_DATA_TEMPR1[71] , 
        \R_DATA_TEMPR2[71] , \R_DATA_TEMPR3[71] , \R_DATA_TEMPR4[71] , 
        \R_DATA_TEMPR5[71] , \R_DATA_TEMPR6[71] , \R_DATA_TEMPR7[71] , 
        \R_DATA_TEMPR8[71] , \R_DATA_TEMPR9[71] , \R_DATA_TEMPR10[71] , 
        \R_DATA_TEMPR11[71] , \R_DATA_TEMPR12[71] , 
        \R_DATA_TEMPR13[71] , \R_DATA_TEMPR14[71] , 
        \R_DATA_TEMPR15[71] , \R_DATA_TEMPR0[72] , \R_DATA_TEMPR1[72] , 
        \R_DATA_TEMPR2[72] , \R_DATA_TEMPR3[72] , \R_DATA_TEMPR4[72] , 
        \R_DATA_TEMPR5[72] , \R_DATA_TEMPR6[72] , \R_DATA_TEMPR7[72] , 
        \R_DATA_TEMPR8[72] , \R_DATA_TEMPR9[72] , \R_DATA_TEMPR10[72] , 
        \R_DATA_TEMPR11[72] , \R_DATA_TEMPR12[72] , 
        \R_DATA_TEMPR13[72] , \R_DATA_TEMPR14[72] , 
        \R_DATA_TEMPR15[72] , \R_DATA_TEMPR0[73] , \R_DATA_TEMPR1[73] , 
        \R_DATA_TEMPR2[73] , \R_DATA_TEMPR3[73] , \R_DATA_TEMPR4[73] , 
        \R_DATA_TEMPR5[73] , \R_DATA_TEMPR6[73] , \R_DATA_TEMPR7[73] , 
        \R_DATA_TEMPR8[73] , \R_DATA_TEMPR9[73] , \R_DATA_TEMPR10[73] , 
        \R_DATA_TEMPR11[73] , \R_DATA_TEMPR12[73] , 
        \R_DATA_TEMPR13[73] , \R_DATA_TEMPR14[73] , 
        \R_DATA_TEMPR15[73] , \R_DATA_TEMPR0[74] , \R_DATA_TEMPR1[74] , 
        \R_DATA_TEMPR2[74] , \R_DATA_TEMPR3[74] , \R_DATA_TEMPR4[74] , 
        \R_DATA_TEMPR5[74] , \R_DATA_TEMPR6[74] , \R_DATA_TEMPR7[74] , 
        \R_DATA_TEMPR8[74] , \R_DATA_TEMPR9[74] , \R_DATA_TEMPR10[74] , 
        \R_DATA_TEMPR11[74] , \R_DATA_TEMPR12[74] , 
        \R_DATA_TEMPR13[74] , \R_DATA_TEMPR14[74] , 
        \R_DATA_TEMPR15[74] , \R_DATA_TEMPR0[75] , \R_DATA_TEMPR1[75] , 
        \R_DATA_TEMPR2[75] , \R_DATA_TEMPR3[75] , \R_DATA_TEMPR4[75] , 
        \R_DATA_TEMPR5[75] , \R_DATA_TEMPR6[75] , \R_DATA_TEMPR7[75] , 
        \R_DATA_TEMPR8[75] , \R_DATA_TEMPR9[75] , \R_DATA_TEMPR10[75] , 
        \R_DATA_TEMPR11[75] , \R_DATA_TEMPR12[75] , 
        \R_DATA_TEMPR13[75] , \R_DATA_TEMPR14[75] , 
        \R_DATA_TEMPR15[75] , \R_DATA_TEMPR0[76] , \R_DATA_TEMPR1[76] , 
        \R_DATA_TEMPR2[76] , \R_DATA_TEMPR3[76] , \R_DATA_TEMPR4[76] , 
        \R_DATA_TEMPR5[76] , \R_DATA_TEMPR6[76] , \R_DATA_TEMPR7[76] , 
        \R_DATA_TEMPR8[76] , \R_DATA_TEMPR9[76] , \R_DATA_TEMPR10[76] , 
        \R_DATA_TEMPR11[76] , \R_DATA_TEMPR12[76] , 
        \R_DATA_TEMPR13[76] , \R_DATA_TEMPR14[76] , 
        \R_DATA_TEMPR15[76] , \R_DATA_TEMPR0[77] , \R_DATA_TEMPR1[77] , 
        \R_DATA_TEMPR2[77] , \R_DATA_TEMPR3[77] , \R_DATA_TEMPR4[77] , 
        \R_DATA_TEMPR5[77] , \R_DATA_TEMPR6[77] , \R_DATA_TEMPR7[77] , 
        \R_DATA_TEMPR8[77] , \R_DATA_TEMPR9[77] , \R_DATA_TEMPR10[77] , 
        \R_DATA_TEMPR11[77] , \R_DATA_TEMPR12[77] , 
        \R_DATA_TEMPR13[77] , \R_DATA_TEMPR14[77] , 
        \R_DATA_TEMPR15[77] , \R_DATA_TEMPR0[78] , \R_DATA_TEMPR1[78] , 
        \R_DATA_TEMPR2[78] , \R_DATA_TEMPR3[78] , \R_DATA_TEMPR4[78] , 
        \R_DATA_TEMPR5[78] , \R_DATA_TEMPR6[78] , \R_DATA_TEMPR7[78] , 
        \R_DATA_TEMPR8[78] , \R_DATA_TEMPR9[78] , \R_DATA_TEMPR10[78] , 
        \R_DATA_TEMPR11[78] , \R_DATA_TEMPR12[78] , 
        \R_DATA_TEMPR13[78] , \R_DATA_TEMPR14[78] , 
        \R_DATA_TEMPR15[78] , \R_DATA_TEMPR0[79] , \R_DATA_TEMPR1[79] , 
        \R_DATA_TEMPR2[79] , \R_DATA_TEMPR3[79] , \R_DATA_TEMPR4[79] , 
        \R_DATA_TEMPR5[79] , \R_DATA_TEMPR6[79] , \R_DATA_TEMPR7[79] , 
        \R_DATA_TEMPR8[79] , \R_DATA_TEMPR9[79] , \R_DATA_TEMPR10[79] , 
        \R_DATA_TEMPR11[79] , \R_DATA_TEMPR12[79] , 
        \R_DATA_TEMPR13[79] , \R_DATA_TEMPR14[79] , 
        \R_DATA_TEMPR15[79] , \BLKX0[0] , \BLKY0[0] , \BLKX1[0] , 
        \BLKY1[0] , \BLKX2[0] , \BLKX2[1] , \BLKX2[2] , \BLKX2[3] , 
        \BLKY2[0] , \BLKY2[1] , \BLKY2[2] , \BLKY2[3] , 
        \ACCESS_BUSY[0][0] , \ACCESS_BUSY[0][1] , \ACCESS_BUSY[1][0] , 
        \ACCESS_BUSY[1][1] , \ACCESS_BUSY[2][0] , \ACCESS_BUSY[2][1] , 
        \ACCESS_BUSY[3][0] , \ACCESS_BUSY[3][1] , \ACCESS_BUSY[4][0] , 
        \ACCESS_BUSY[4][1] , \ACCESS_BUSY[5][0] , \ACCESS_BUSY[5][1] , 
        \ACCESS_BUSY[6][0] , \ACCESS_BUSY[6][1] , \ACCESS_BUSY[7][0] , 
        \ACCESS_BUSY[7][1] , \ACCESS_BUSY[8][0] , \ACCESS_BUSY[8][1] , 
        \ACCESS_BUSY[9][0] , \ACCESS_BUSY[9][1] , \ACCESS_BUSY[10][0] , 
        \ACCESS_BUSY[10][1] , \ACCESS_BUSY[11][0] , 
        \ACCESS_BUSY[11][1] , \ACCESS_BUSY[12][0] , 
        \ACCESS_BUSY[12][1] , \ACCESS_BUSY[13][0] , 
        \ACCESS_BUSY[13][1] , \ACCESS_BUSY[14][0] , 
        \ACCESS_BUSY[14][1] , \ACCESS_BUSY[15][0] , 
        \ACCESS_BUSY[15][1] , OR4_31_Y, OR4_203_Y, OR4_5_Y, OR4_262_Y, 
        OR4_265_Y, OR4_68_Y, OR4_306_Y, OR4_84_Y, OR4_217_Y, OR4_174_Y, 
        OR4_78_Y, OR4_108_Y, OR4_239_Y, OR4_162_Y, OR4_76_Y, OR4_12_Y, 
        OR4_314_Y, OR4_288_Y, OR4_188_Y, OR4_222_Y, OR4_137_Y, 
        OR4_126_Y, OR4_273_Y, OR4_245_Y, OR4_92_Y, OR4_299_Y, 
        OR4_124_Y, OR4_234_Y, OR4_20_Y, OR4_98_Y, OR4_50_Y, OR4_79_Y, 
        OR4_266_Y, OR4_69_Y, OR4_307_Y, OR4_85_Y, OR4_210_Y, OR4_91_Y, 
        OR4_232_Y, OR4_24_Y, OR4_105_Y, OR4_176_Y, OR4_130_Y, 
        OR4_152_Y, OR4_315_Y, OR4_224_Y, OR4_144_Y, OR4_298_Y, 
        OR4_106_Y, OR4_177_Y, OR4_131_Y, OR4_153_Y, OR4_276_Y, 
        OR4_88_Y, OR4_291_Y, OR4_237_Y, OR4_235_Y, OR4_75_Y, OR4_213_Y, 
        OR4_142_Y, OR4_13_Y, OR4_2_Y, OR4_148_Y, OR4_123_Y, OR4_145_Y, 
        OR4_264_Y, OR4_184_Y, OR4_283_Y, OR4_280_Y, OR4_115_Y, 
        OR4_250_Y, OR4_183_Y, OR4_209_Y, OR4_166_Y, OR4_70_Y, 
        OR4_104_Y, OR4_77_Y, OR4_229_Y, OR4_32_Y, OR4_295_Y, OR4_63_Y, 
        OR4_18_Y, OR4_253_Y, OR4_111_Y, OR4_211_Y, OR4_287_Y, 
        OR4_180_Y, OR4_94_Y, OR4_64_Y, OR4_45_Y, OR4_202_Y, OR4_161_Y, 
        OR4_194_Y, OR4_310_Y, OR4_228_Y, OR4_6_Y, OR4_46_Y, OR4_305_Y, 
        OR4_221_Y, OR4_218_Y, OR4_86_Y, OR4_293_Y, OR4_116_Y, 
        OR4_230_Y, OR4_167_Y, OR4_156_Y, OR4_308_Y, OR4_275_Y, 
        OR4_301_Y, OR4_101_Y, OR4_16_Y, OR4_119_Y, OR4_267_Y, OR4_57_Y, 
        OR4_196_Y, OR4_34_Y, OR4_128_Y, OR4_268_Y, OR4_117_Y, 
        OR4_289_Y, OR4_138_Y, OR4_102_Y, OR4_8_Y, OR4_195_Y, OR4_279_Y, 
        OR4_38_Y, OR4_259_Y, OR4_171_Y, OR4_302_Y, OR4_58_Y, OR4_7_Y, 
        OR4_27_Y, OR4_139_Y, OR4_103_Y, OR4_9_Y, OR4_197_Y, OR4_281_Y, 
        OR4_39_Y, OR4_261_Y, OR4_172_Y, OR4_22_Y, OR4_132_Y, OR4_269_Y, 
        OR4_120_Y, OR4_21_Y, OR4_100_Y, OR4_54_Y, OR4_80_Y, OR4_140_Y, 
        OR4_220_Y, OR4_159_Y, OR4_190_Y, OR4_23_Y, OR4_133_Y, 
        OR4_271_Y, OR4_121_Y, OR4_274_Y, OR4_110_Y, OR4_243_Y, 
        OR4_179_Y, OR4_41_Y, OR4_236_Y, OR4_146_Y, OR4_134_Y, OR4_55_Y, 
        OR4_37_Y, OR4_193_Y, OR4_157_Y, OR4_187_Y, OR4_303_Y, 
        OR4_223_Y, OR4_319_Y, OR4_25_Y, OR4_241_Y, OR4_231_Y, OR4_53_Y, 
        OR4_14_Y, OR4_300_Y, OR4_219_Y, OR4_71_Y, OR4_155_Y, OR4_240_Y, 
        OR4_141_Y, OR4_48_Y, OR4_118_Y, OR4_143_Y, OR4_74_Y, OR4_204_Y, 
        OR4_282_Y, OR4_93_Y, OR4_292_Y, OR4_242_Y, OR4_226_Y, OR4_11_Y, 
        OR4_147_Y, OR4_316_Y, OR4_65_Y, OR4_19_Y, OR4_255_Y, OR4_112_Y, 
        OR4_212_Y, OR4_290_Y, OR4_182_Y, OR4_97_Y, OR4_170_Y, 
        OR4_135_Y, OR4_40_Y, OR4_225_Y, OR4_313_Y, OR4_82_Y, OR4_294_Y, 
        OR4_216_Y, OR4_17_Y, OR4_96_Y, OR4_44_Y, OR4_72_Y, OR4_270_Y, 
        OR4_60_Y, OR4_198_Y, OR4_36_Y, OR4_215_Y, OR4_173_Y, OR4_73_Y, 
        OR4_107_Y, OR4_66_Y, OR4_163_Y, OR4_304_Y, OR4_154_Y, 
        OR4_114_Y, OR4_256_Y, OR4_175_Y, OR4_10_Y, OR4_33_Y, OR4_168_Y, 
        OR4_51_Y, OR4_317_Y, OR4_90_Y, OR4_297_Y, OR4_122_Y, OR4_233_Y, 
        OR4_35_Y, OR4_169_Y, OR4_52_Y, OR4_318_Y, OR4_284_Y, OR4_252_Y, 
        OR4_149_Y, OR4_185_Y, OR4_164_Y, OR4_59_Y, OR4_206_Y, 
        OR4_311_Y, OR4_286_Y, OR4_254_Y, OR4_151_Y, OR4_186_Y, 
        OR4_165_Y, OR4_61_Y, OR4_207_Y, OR4_312_Y, OR4_56_Y, OR4_15_Y, 
        OR4_249_Y, OR4_109_Y, OR4_205_Y, OR4_278_Y, OR4_178_Y, 
        OR4_89_Y, OR4_277_Y, OR4_113_Y, OR4_248_Y, OR4_181_Y, 
        OR4_258_Y, OR4_0_Y, OR4_191_Y, OR4_99_Y, OR4_263_Y, OR4_49_Y, 
        OR4_189_Y, OR4_29_Y, OR4_238_Y, OR4_47_Y, OR4_251_Y, OR4_208_Y, 
        OR4_62_Y, OR4_43_Y, OR4_199_Y, OR4_160_Y, OR4_192_Y, OR4_309_Y, 
        OR4_227_Y, OR4_4_Y, OR4_285_Y, OR4_95_Y, OR4_296_Y, OR4_246_Y, 
        OR4_247_Y, OR4_127_Y, OR4_150_Y, OR4_1_Y, OR4_158_Y, OR4_129_Y, 
        OR4_26_Y, OR4_67_Y, OR4_81_Y, OR4_214_Y, OR4_87_Y, OR4_28_Y, 
        OR4_30_Y, OR4_201_Y, OR4_3_Y, OR4_260_Y, OR4_42_Y, OR4_257_Y, 
        OR4_83_Y, OR4_200_Y, OR4_136_Y, OR4_125_Y, OR4_272_Y, 
        OR4_244_Y, VCC, GND, ADLIB_VCC;
    wire GND_power_net1;
    wire VCC_power_net1;
    assign GND = GND_power_net1;
    assign VCC = VCC_power_net1;
    assign ADLIB_VCC = VCC_power_net1;
    
    OR4 OR4_172 (.A(\R_DATA_TEMPR12[78] ), .B(\R_DATA_TEMPR13[78] ), 
        .C(\R_DATA_TEMPR14[78] ), .D(\R_DATA_TEMPR15[78] ), .Y(
        OR4_172_Y));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%9%1%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C1 (.A_DOUT({
        \R_DATA_TEMPR9[79] , \R_DATA_TEMPR9[78] , \R_DATA_TEMPR9[77] , 
        \R_DATA_TEMPR9[76] , \R_DATA_TEMPR9[75] , \R_DATA_TEMPR9[74] , 
        \R_DATA_TEMPR9[73] , \R_DATA_TEMPR9[72] , \R_DATA_TEMPR9[71] , 
        \R_DATA_TEMPR9[70] , \R_DATA_TEMPR9[69] , \R_DATA_TEMPR9[68] , 
        \R_DATA_TEMPR9[67] , \R_DATA_TEMPR9[66] , \R_DATA_TEMPR9[65] , 
        \R_DATA_TEMPR9[64] , \R_DATA_TEMPR9[63] , \R_DATA_TEMPR9[62] , 
        \R_DATA_TEMPR9[61] , \R_DATA_TEMPR9[60] }), .B_DOUT({
        \R_DATA_TEMPR9[59] , \R_DATA_TEMPR9[58] , \R_DATA_TEMPR9[57] , 
        \R_DATA_TEMPR9[56] , \R_DATA_TEMPR9[55] , \R_DATA_TEMPR9[54] , 
        \R_DATA_TEMPR9[53] , \R_DATA_TEMPR9[52] , \R_DATA_TEMPR9[51] , 
        \R_DATA_TEMPR9[50] , \R_DATA_TEMPR9[49] , \R_DATA_TEMPR9[48] , 
        \R_DATA_TEMPR9[47] , \R_DATA_TEMPR9[46] , \R_DATA_TEMPR9[45] , 
        \R_DATA_TEMPR9[44] , \R_DATA_TEMPR9[43] , \R_DATA_TEMPR9[42] , 
        \R_DATA_TEMPR9[41] , \R_DATA_TEMPR9[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[9][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[2] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_145 (.A(\R_DATA_TEMPR0[54] ), .B(\R_DATA_TEMPR1[54] ), .C(
        \R_DATA_TEMPR2[54] ), .D(\R_DATA_TEMPR3[54] ), .Y(OR4_145_Y));
    OR4 OR4_31 (.A(\R_DATA_TEMPR0[73] ), .B(\R_DATA_TEMPR1[73] ), .C(
        \R_DATA_TEMPR2[73] ), .D(\R_DATA_TEMPR3[73] ), .Y(OR4_31_Y));
    OR4 \OR4_R_DATA[21]  (.A(OR4_217_Y), .B(OR4_174_Y), .C(OR4_78_Y), 
        .D(OR4_108_Y), .Y(R_DATA[21]));
    OR4 \OR4_R_DATA[37]  (.A(OR4_33_Y), .B(OR4_168_Y), .C(OR4_51_Y), 
        .D(OR4_317_Y), .Y(R_DATA[37]));
    OR4 OR4_296 (.A(\R_DATA_TEMPR8[27] ), .B(\R_DATA_TEMPR9[27] ), .C(
        \R_DATA_TEMPR10[27] ), .D(\R_DATA_TEMPR11[27] ), .Y(OR4_296_Y));
    OR4 OR4_14 (.A(\R_DATA_TEMPR0[59] ), .B(\R_DATA_TEMPR1[59] ), .C(
        \R_DATA_TEMPR2[59] ), .D(\R_DATA_TEMPR3[59] ), .Y(OR4_14_Y));
    OR4 OR4_64 (.A(\R_DATA_TEMPR0[25] ), .B(\R_DATA_TEMPR1[25] ), .C(
        \R_DATA_TEMPR2[25] ), .D(\R_DATA_TEMPR3[25] ), .Y(OR4_64_Y));
    OR4 \OR4_R_DATA[59]  (.A(OR4_14_Y), .B(OR4_300_Y), .C(OR4_219_Y), 
        .D(OR4_71_Y), .Y(R_DATA[59]));
    OR4 OR4_194 (.A(\R_DATA_TEMPR0[24] ), .B(\R_DATA_TEMPR1[24] ), .C(
        \R_DATA_TEMPR2[24] ), .D(\R_DATA_TEMPR3[24] ), .Y(OR4_194_Y));
    OR4 OR4_108 (.A(\R_DATA_TEMPR12[21] ), .B(\R_DATA_TEMPR13[21] ), 
        .C(\R_DATA_TEMPR14[21] ), .D(\R_DATA_TEMPR15[21] ), .Y(
        OR4_108_Y));
    OR4 \OR4_R_DATA[17]  (.A(OR4_282_Y), .B(OR4_93_Y), .C(OR4_292_Y), 
        .D(OR4_242_Y), .Y(R_DATA[17]));
    OR4 OR4_293 (.A(\R_DATA_TEMPR4[62] ), .B(\R_DATA_TEMPR5[62] ), .C(
        \R_DATA_TEMPR6[62] ), .D(\R_DATA_TEMPR7[62] ), .Y(OR4_293_Y));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%5%0%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C0 (.A_DOUT({
        \R_DATA_TEMPR5[39] , \R_DATA_TEMPR5[38] , \R_DATA_TEMPR5[37] , 
        \R_DATA_TEMPR5[36] , \R_DATA_TEMPR5[35] , \R_DATA_TEMPR5[34] , 
        \R_DATA_TEMPR5[33] , \R_DATA_TEMPR5[32] , \R_DATA_TEMPR5[31] , 
        \R_DATA_TEMPR5[30] , \R_DATA_TEMPR5[29] , \R_DATA_TEMPR5[28] , 
        \R_DATA_TEMPR5[27] , \R_DATA_TEMPR5[26] , \R_DATA_TEMPR5[25] , 
        \R_DATA_TEMPR5[24] , \R_DATA_TEMPR5[23] , \R_DATA_TEMPR5[22] , 
        \R_DATA_TEMPR5[21] , \R_DATA_TEMPR5[20] }), .B_DOUT({
        \R_DATA_TEMPR5[19] , \R_DATA_TEMPR5[18] , \R_DATA_TEMPR5[17] , 
        \R_DATA_TEMPR5[16] , \R_DATA_TEMPR5[15] , \R_DATA_TEMPR5[14] , 
        \R_DATA_TEMPR5[13] , \R_DATA_TEMPR5[12] , \R_DATA_TEMPR5[11] , 
        \R_DATA_TEMPR5[10] , \R_DATA_TEMPR5[9] , \R_DATA_TEMPR5[8] , 
        \R_DATA_TEMPR5[7] , \R_DATA_TEMPR5[6] , \R_DATA_TEMPR5[5] , 
        \R_DATA_TEMPR5[4] , \R_DATA_TEMPR5[3] , \R_DATA_TEMPR5[2] , 
        \R_DATA_TEMPR5[1] , \R_DATA_TEMPR5[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[5][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[1] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_261 (.A(\R_DATA_TEMPR8[78] ), .B(\R_DATA_TEMPR9[78] ), .C(
        \R_DATA_TEMPR10[78] ), .D(\R_DATA_TEMPR11[78] ), .Y(OR4_261_Y));
    OR4 OR4_312 (.A(\R_DATA_TEMPR12[72] ), .B(\R_DATA_TEMPR13[72] ), 
        .C(\R_DATA_TEMPR14[72] ), .D(\R_DATA_TEMPR15[72] ), .Y(
        OR4_312_Y));
    OR4 OR4_249 (.A(\R_DATA_TEMPR8[69] ), .B(\R_DATA_TEMPR9[69] ), .C(
        \R_DATA_TEMPR10[69] ), .D(\R_DATA_TEMPR11[69] ), .Y(OR4_249_Y));
    OR4 \OR4_R_DATA[3]  (.A(OR4_128_Y), .B(OR4_268_Y), .C(OR4_117_Y), 
        .D(OR4_289_Y), .Y(R_DATA[3]));
    OR4 OR4_109 (.A(\R_DATA_TEMPR12[69] ), .B(\R_DATA_TEMPR13[69] ), 
        .C(\R_DATA_TEMPR14[69] ), .D(\R_DATA_TEMPR15[69] ), .Y(
        OR4_109_Y));
    OR4 OR4_56 (.A(\R_DATA_TEMPR0[69] ), .B(\R_DATA_TEMPR1[69] ), .C(
        \R_DATA_TEMPR2[69] ), .D(\R_DATA_TEMPR3[69] ), .Y(OR4_56_Y));
    OR4 OR4_294 (.A(\R_DATA_TEMPR8[48] ), .B(\R_DATA_TEMPR9[48] ), .C(
        \R_DATA_TEMPR10[48] ), .D(\R_DATA_TEMPR11[48] ), .Y(OR4_294_Y));
    OR4 OR4_123 (.A(\R_DATA_TEMPR12[55] ), .B(\R_DATA_TEMPR13[55] ), 
        .C(\R_DATA_TEMPR14[55] ), .D(\R_DATA_TEMPR15[55] ), .Y(
        OR4_123_Y));
    OR4 OR4_96 (.A(\R_DATA_TEMPR4[66] ), .B(\R_DATA_TEMPR5[66] ), .C(
        \R_DATA_TEMPR6[66] ), .D(\R_DATA_TEMPR7[66] ), .Y(OR4_96_Y));
    CFG3 #( .INIT(8'h20) )  \CFG3_BLKX2[2]  (.A(W_ADDR[12]), .B(
        W_ADDR[11]), .C(W_EN), .Y(\BLKX2[2] ));
    OR4 OR4_105 (.A(\R_DATA_TEMPR0[36] ), .B(\R_DATA_TEMPR1[36] ), .C(
        \R_DATA_TEMPR2[36] ), .D(\R_DATA_TEMPR3[36] ), .Y(OR4_105_Y));
    OR4 \OR4_R_DATA[48]  (.A(OR4_313_Y), .B(OR4_82_Y), .C(OR4_294_Y), 
        .D(OR4_216_Y), .Y(R_DATA[48]));
    OR4 OR4_0 (.A(\R_DATA_TEMPR4[7] ), .B(\R_DATA_TEMPR5[7] ), .C(
        \R_DATA_TEMPR6[7] ), .D(\R_DATA_TEMPR7[7] ), .Y(OR4_0_Y));
    OR4 \OR4_R_DATA[46]  (.A(OR4_140_Y), .B(OR4_220_Y), .C(OR4_159_Y), 
        .D(OR4_190_Y), .Y(R_DATA[46]));
    OR4 OR4_131 (.A(\R_DATA_TEMPR8[76] ), .B(\R_DATA_TEMPR9[76] ), .C(
        \R_DATA_TEMPR10[76] ), .D(\R_DATA_TEMPR11[76] ), .Y(OR4_131_Y));
    OR4 OR4_197 (.A(\R_DATA_TEMPR12[79] ), .B(\R_DATA_TEMPR13[79] ), 
        .C(\R_DATA_TEMPR14[79] ), .D(\R_DATA_TEMPR15[79] ), .Y(
        OR4_197_Y));
    OR4 OR4_10 (.A(\R_DATA_TEMPR12[5] ), .B(\R_DATA_TEMPR13[5] ), .C(
        \R_DATA_TEMPR14[5] ), .D(\R_DATA_TEMPR15[5] ), .Y(OR4_10_Y));
    OR4 OR4_60 (.A(\R_DATA_TEMPR4[20] ), .B(\R_DATA_TEMPR5[20] ), .C(
        \R_DATA_TEMPR6[20] ), .D(\R_DATA_TEMPR7[20] ), .Y(OR4_60_Y));
    OR4 \OR4_R_DATA[30]  (.A(OR4_22_Y), .B(OR4_132_Y), .C(OR4_269_Y), 
        .D(OR4_120_Y), .Y(R_DATA[30]));
    OR4 OR4_173 (.A(\R_DATA_TEMPR4[11] ), .B(\R_DATA_TEMPR5[11] ), .C(
        \R_DATA_TEMPR6[11] ), .D(\R_DATA_TEMPR7[11] ), .Y(OR4_173_Y));
    OR4 OR4_255 (.A(\R_DATA_TEMPR8[29] ), .B(\R_DATA_TEMPR9[29] ), .C(
        \R_DATA_TEMPR10[29] ), .D(\R_DATA_TEMPR11[29] ), .Y(OR4_255_Y));
    OR4 OR4_25 (.A(\R_DATA_TEMPR0[2] ), .B(\R_DATA_TEMPR1[2] ), .C(
        \R_DATA_TEMPR2[2] ), .D(\R_DATA_TEMPR3[2] ), .Y(OR4_25_Y));
    OR4 \OR4_R_DATA[10]  (.A(OR4_267_Y), .B(OR4_57_Y), .C(OR4_196_Y), 
        .D(OR4_34_Y), .Y(R_DATA[10]));
    OR4 OR4_209 (.A(\R_DATA_TEMPR0[61] ), .B(\R_DATA_TEMPR1[61] ), .C(
        \R_DATA_TEMPR2[61] ), .D(\R_DATA_TEMPR3[61] ), .Y(OR4_209_Y));
    OR4 OR4_215 (.A(\R_DATA_TEMPR0[11] ), .B(\R_DATA_TEMPR1[11] ), .C(
        \R_DATA_TEMPR2[11] ), .D(\R_DATA_TEMPR3[11] ), .Y(OR4_215_Y));
    OR4 OR4_21 (.A(\R_DATA_TEMPR0[26] ), .B(\R_DATA_TEMPR1[26] ), .C(
        \R_DATA_TEMPR2[26] ), .D(\R_DATA_TEMPR3[26] ), .Y(OR4_21_Y));
    OR4 \OR4_R_DATA[24]  (.A(OR4_194_Y), .B(OR4_310_Y), .C(OR4_228_Y), 
        .D(OR4_6_Y), .Y(R_DATA[24]));
    OR4 OR4_89 (.A(\R_DATA_TEMPR12[68] ), .B(\R_DATA_TEMPR13[68] ), .C(
        \R_DATA_TEMPR14[68] ), .D(\R_DATA_TEMPR15[68] ), .Y(OR4_89_Y));
    OR4 OR4_287 (.A(\R_DATA_TEMPR4[18] ), .B(\R_DATA_TEMPR5[18] ), .C(
        \R_DATA_TEMPR6[18] ), .D(\R_DATA_TEMPR7[18] ), .Y(OR4_287_Y));
    OR4 \OR4_R_DATA[23]  (.A(OR4_280_Y), .B(OR4_115_Y), .C(OR4_250_Y), 
        .D(OR4_183_Y), .Y(R_DATA[23]));
    OR4 OR4_250 (.A(\R_DATA_TEMPR8[23] ), .B(\R_DATA_TEMPR9[23] ), .C(
        \R_DATA_TEMPR10[23] ), .D(\R_DATA_TEMPR11[23] ), .Y(OR4_250_Y));
    OR4 OR4_46 (.A(\R_DATA_TEMPR0[9] ), .B(\R_DATA_TEMPR1[9] ), .C(
        \R_DATA_TEMPR2[9] ), .D(\R_DATA_TEMPR3[9] ), .Y(OR4_46_Y));
    OR4 OR4_138 (.A(\R_DATA_TEMPR0[39] ), .B(\R_DATA_TEMPR1[39] ), .C(
        \R_DATA_TEMPR2[39] ), .D(\R_DATA_TEMPR3[39] ), .Y(OR4_138_Y));
    OR4 OR4_298 (.A(\R_DATA_TEMPR12[0] ), .B(\R_DATA_TEMPR13[0] ), .C(
        \R_DATA_TEMPR14[0] ), .D(\R_DATA_TEMPR15[0] ), .Y(OR4_298_Y));
    OR4 \OR4_R_DATA[57]  (.A(OR4_238_Y), .B(OR4_47_Y), .C(OR4_251_Y), 
        .D(OR4_208_Y), .Y(R_DATA[57]));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%5%1%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C1 (.A_DOUT({
        \R_DATA_TEMPR5[79] , \R_DATA_TEMPR5[78] , \R_DATA_TEMPR5[77] , 
        \R_DATA_TEMPR5[76] , \R_DATA_TEMPR5[75] , \R_DATA_TEMPR5[74] , 
        \R_DATA_TEMPR5[73] , \R_DATA_TEMPR5[72] , \R_DATA_TEMPR5[71] , 
        \R_DATA_TEMPR5[70] , \R_DATA_TEMPR5[69] , \R_DATA_TEMPR5[68] , 
        \R_DATA_TEMPR5[67] , \R_DATA_TEMPR5[66] , \R_DATA_TEMPR5[65] , 
        \R_DATA_TEMPR5[64] , \R_DATA_TEMPR5[63] , \R_DATA_TEMPR5[62] , 
        \R_DATA_TEMPR5[61] , \R_DATA_TEMPR5[60] }), .B_DOUT({
        \R_DATA_TEMPR5[59] , \R_DATA_TEMPR5[58] , \R_DATA_TEMPR5[57] , 
        \R_DATA_TEMPR5[56] , \R_DATA_TEMPR5[55] , \R_DATA_TEMPR5[54] , 
        \R_DATA_TEMPR5[53] , \R_DATA_TEMPR5[52] , \R_DATA_TEMPR5[51] , 
        \R_DATA_TEMPR5[50] , \R_DATA_TEMPR5[49] , \R_DATA_TEMPR5[48] , 
        \R_DATA_TEMPR5[47] , \R_DATA_TEMPR5[46] , \R_DATA_TEMPR5[45] , 
        \R_DATA_TEMPR5[44] , \R_DATA_TEMPR5[43] , \R_DATA_TEMPR5[42] , 
        \R_DATA_TEMPR5[41] , \R_DATA_TEMPR5[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[5][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[1] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_246 (.A(\R_DATA_TEMPR12[27] ), .B(\R_DATA_TEMPR13[27] ), 
        .C(\R_DATA_TEMPR14[27] ), .D(\R_DATA_TEMPR15[27] ), .Y(
        OR4_246_Y));
    OR4 OR4_210 (.A(\R_DATA_TEMPR0[42] ), .B(\R_DATA_TEMPR1[42] ), .C(
        \R_DATA_TEMPR2[42] ), .D(\R_DATA_TEMPR3[42] ), .Y(OR4_210_Y));
    OR4 OR4_144 (.A(\R_DATA_TEMPR8[0] ), .B(\R_DATA_TEMPR9[0] ), .C(
        \R_DATA_TEMPR10[0] ), .D(\R_DATA_TEMPR11[0] ), .Y(OR4_144_Y));
    OR4 \OR4_R_DATA[25]  (.A(OR4_64_Y), .B(OR4_45_Y), .C(OR4_202_Y), 
        .D(OR4_161_Y), .Y(R_DATA[25]));
    OR4 OR4_243 (.A(\R_DATA_TEMPR8[63] ), .B(\R_DATA_TEMPR9[63] ), .C(
        \R_DATA_TEMPR10[63] ), .D(\R_DATA_TEMPR11[63] ), .Y(OR4_243_Y));
    OR4 OR4_221 (.A(\R_DATA_TEMPR8[9] ), .B(\R_DATA_TEMPR9[9] ), .C(
        \R_DATA_TEMPR10[9] ), .D(\R_DATA_TEMPR11[9] ), .Y(OR4_221_Y));
    OR4 OR4_139 (.A(\R_DATA_TEMPR0[79] ), .B(\R_DATA_TEMPR1[79] ), .C(
        \R_DATA_TEMPR2[79] ), .D(\R_DATA_TEMPR3[79] ), .Y(OR4_139_Y));
    OR4 \OR4_R_DATA[7]  (.A(OR4_258_Y), .B(OR4_0_Y), .C(OR4_191_Y), .D(
        OR4_99_Y), .Y(R_DATA[7]));
    OR4 OR4_52 (.A(\R_DATA_TEMPR8[77] ), .B(\R_DATA_TEMPR9[77] ), .C(
        \R_DATA_TEMPR10[77] ), .D(\R_DATA_TEMPR11[77] ), .Y(OR4_52_Y));
    OR4 OR4_92 (.A(\R_DATA_TEMPR0[22] ), .B(\R_DATA_TEMPR1[22] ), .C(
        \R_DATA_TEMPR2[22] ), .D(\R_DATA_TEMPR3[22] ), .Y(OR4_92_Y));
    OR4 OR4_244 (.A(\R_DATA_TEMPR12[35] ), .B(\R_DATA_TEMPR13[35] ), 
        .C(\R_DATA_TEMPR14[35] ), .D(\R_DATA_TEMPR15[35] ), .Y(
        OR4_244_Y));
    OR4 OR4_79 (.A(\R_DATA_TEMPR12[16] ), .B(\R_DATA_TEMPR13[16] ), .C(
        \R_DATA_TEMPR14[16] ), .D(\R_DATA_TEMPR15[16] ), .Y(OR4_79_Y));
    OR4 OR4_135 (.A(\R_DATA_TEMPR4[49] ), .B(\R_DATA_TEMPR5[49] ), .C(
        \R_DATA_TEMPR6[49] ), .D(\R_DATA_TEMPR7[49] ), .Y(OR4_135_Y));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%14%0%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C0 (.A_DOUT({
        \R_DATA_TEMPR14[39] , \R_DATA_TEMPR14[38] , 
        \R_DATA_TEMPR14[37] , \R_DATA_TEMPR14[36] , 
        \R_DATA_TEMPR14[35] , \R_DATA_TEMPR14[34] , 
        \R_DATA_TEMPR14[33] , \R_DATA_TEMPR14[32] , 
        \R_DATA_TEMPR14[31] , \R_DATA_TEMPR14[30] , 
        \R_DATA_TEMPR14[29] , \R_DATA_TEMPR14[28] , 
        \R_DATA_TEMPR14[27] , \R_DATA_TEMPR14[26] , 
        \R_DATA_TEMPR14[25] , \R_DATA_TEMPR14[24] , 
        \R_DATA_TEMPR14[23] , \R_DATA_TEMPR14[22] , 
        \R_DATA_TEMPR14[21] , \R_DATA_TEMPR14[20] }), .B_DOUT({
        \R_DATA_TEMPR14[19] , \R_DATA_TEMPR14[18] , 
        \R_DATA_TEMPR14[17] , \R_DATA_TEMPR14[16] , 
        \R_DATA_TEMPR14[15] , \R_DATA_TEMPR14[14] , 
        \R_DATA_TEMPR14[13] , \R_DATA_TEMPR14[12] , 
        \R_DATA_TEMPR14[11] , \R_DATA_TEMPR14[10] , 
        \R_DATA_TEMPR14[9] , \R_DATA_TEMPR14[8] , \R_DATA_TEMPR14[7] , 
        \R_DATA_TEMPR14[6] , \R_DATA_TEMPR14[5] , \R_DATA_TEMPR14[4] , 
        \R_DATA_TEMPR14[3] , \R_DATA_TEMPR14[2] , \R_DATA_TEMPR14[1] , 
        \R_DATA_TEMPR14[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[14][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[3] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[3] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_252 (.A(\R_DATA_TEMPR4[31] ), .B(\R_DATA_TEMPR5[31] ), .C(
        \R_DATA_TEMPR6[31] ), .D(\R_DATA_TEMPR7[31] ), .Y(OR4_252_Y));
    OR4 OR4_271 (.A(\R_DATA_TEMPR8[70] ), .B(\R_DATA_TEMPR9[70] ), .C(
        \R_DATA_TEMPR10[70] ), .D(\R_DATA_TEMPR11[70] ), .Y(OR4_271_Y));
    OR4 OR4_307 (.A(\R_DATA_TEMPR8[74] ), .B(\R_DATA_TEMPR9[74] ), .C(
        \R_DATA_TEMPR10[74] ), .D(\R_DATA_TEMPR11[74] ), .Y(OR4_307_Y));
    OR4 OR4_63 (.A(\R_DATA_TEMPR0[19] ), .B(\R_DATA_TEMPR1[19] ), .C(
        \R_DATA_TEMPR2[19] ), .D(\R_DATA_TEMPR3[19] ), .Y(OR4_63_Y));
    OR4 OR4_13 (.A(\R_DATA_TEMPR0[55] ), .B(\R_DATA_TEMPR1[55] ), .C(
        \R_DATA_TEMPR2[55] ), .D(\R_DATA_TEMPR3[55] ), .Y(OR4_13_Y));
    OR4 OR4_152 (.A(\R_DATA_TEMPR12[36] ), .B(\R_DATA_TEMPR13[36] ), 
        .C(\R_DATA_TEMPR14[36] ), .D(\R_DATA_TEMPR15[36] ), .Y(
        OR4_152_Y));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%9%0%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C0 (.A_DOUT({
        \R_DATA_TEMPR9[39] , \R_DATA_TEMPR9[38] , \R_DATA_TEMPR9[37] , 
        \R_DATA_TEMPR9[36] , \R_DATA_TEMPR9[35] , \R_DATA_TEMPR9[34] , 
        \R_DATA_TEMPR9[33] , \R_DATA_TEMPR9[32] , \R_DATA_TEMPR9[31] , 
        \R_DATA_TEMPR9[30] , \R_DATA_TEMPR9[29] , \R_DATA_TEMPR9[28] , 
        \R_DATA_TEMPR9[27] , \R_DATA_TEMPR9[26] , \R_DATA_TEMPR9[25] , 
        \R_DATA_TEMPR9[24] , \R_DATA_TEMPR9[23] , \R_DATA_TEMPR9[22] , 
        \R_DATA_TEMPR9[21] , \R_DATA_TEMPR9[20] }), .B_DOUT({
        \R_DATA_TEMPR9[19] , \R_DATA_TEMPR9[18] , \R_DATA_TEMPR9[17] , 
        \R_DATA_TEMPR9[16] , \R_DATA_TEMPR9[15] , \R_DATA_TEMPR9[14] , 
        \R_DATA_TEMPR9[13] , \R_DATA_TEMPR9[12] , \R_DATA_TEMPR9[11] , 
        \R_DATA_TEMPR9[10] , \R_DATA_TEMPR9[9] , \R_DATA_TEMPR9[8] , 
        \R_DATA_TEMPR9[7] , \R_DATA_TEMPR9[6] , \R_DATA_TEMPR9[5] , 
        \R_DATA_TEMPR9[4] , \R_DATA_TEMPR9[3] , \R_DATA_TEMPR9[2] , 
        \R_DATA_TEMPR9[1] , \R_DATA_TEMPR9[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[9][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[2] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_57 (.A(\R_DATA_TEMPR4[10] ), .B(\R_DATA_TEMPR5[10] ), .C(
        \R_DATA_TEMPR6[10] ), .D(\R_DATA_TEMPR7[10] ), .Y(OR4_57_Y));
    OR4 OR4_97 (.A(\R_DATA_TEMPR12[28] ), .B(\R_DATA_TEMPR13[28] ), .C(
        \R_DATA_TEMPR14[28] ), .D(\R_DATA_TEMPR15[28] ), .Y(OR4_97_Y));
    OR4 OR4_206 (.A(\R_DATA_TEMPR8[32] ), .B(\R_DATA_TEMPR9[32] ), .C(
        \R_DATA_TEMPR10[32] ), .D(\R_DATA_TEMPR11[32] ), .Y(OR4_206_Y));
    OR4 OR4_181 (.A(\R_DATA_TEMPR12[13] ), .B(\R_DATA_TEMPR13[13] ), 
        .C(\R_DATA_TEMPR14[13] ), .D(\R_DATA_TEMPR15[13] ), .Y(
        OR4_181_Y));
    OR4 OR4_147 (.A(\R_DATA_TEMPR8[50] ), .B(\R_DATA_TEMPR9[50] ), .C(
        \R_DATA_TEMPR10[50] ), .D(\R_DATA_TEMPR11[50] ), .Y(OR4_147_Y));
    OR4 OR4_212 (.A(\R_DATA_TEMPR0[28] ), .B(\R_DATA_TEMPR1[28] ), .C(
        \R_DATA_TEMPR2[28] ), .D(\R_DATA_TEMPR3[28] ), .Y(OR4_212_Y));
    OR4 \OR4_R_DATA[50]  (.A(OR4_226_Y), .B(OR4_11_Y), .C(OR4_147_Y), 
        .D(OR4_316_Y), .Y(R_DATA[50]));
    OR4 OR4_104 (.A(\R_DATA_TEMPR12[61] ), .B(\R_DATA_TEMPR13[61] ), 
        .C(\R_DATA_TEMPR14[61] ), .D(\R_DATA_TEMPR15[61] ), .Y(
        OR4_104_Y));
    OR4 \OR4_R_DATA[22]  (.A(OR4_92_Y), .B(OR4_299_Y), .C(OR4_124_Y), 
        .D(OR4_234_Y), .Y(R_DATA[22]));
    OR4 OR4_239 (.A(\R_DATA_TEMPR0[4] ), .B(\R_DATA_TEMPR1[4] ), .C(
        \R_DATA_TEMPR2[4] ), .D(\R_DATA_TEMPR3[4] ), .Y(OR4_239_Y));
    OR4 OR4_1 (.A(\R_DATA_TEMPR12[1] ), .B(\R_DATA_TEMPR13[1] ), .C(
        \R_DATA_TEMPR14[1] ), .D(\R_DATA_TEMPR15[1] ), .Y(OR4_1_Y));
    OR4 OR4_6 (.A(\R_DATA_TEMPR12[24] ), .B(\R_DATA_TEMPR13[24] ), .C(
        \R_DATA_TEMPR14[24] ), .D(\R_DATA_TEMPR15[24] ), .Y(OR4_6_Y));
    CFG3 #( .INIT(8'h10) )  \CFG3_BLKX2[0]  (.A(W_ADDR[12]), .B(
        W_ADDR[11]), .C(W_EN), .Y(\BLKX2[0] ));
    OR4 OR4_203 (.A(\R_DATA_TEMPR4[73] ), .B(\R_DATA_TEMPR5[73] ), .C(
        \R_DATA_TEMPR6[73] ), .D(\R_DATA_TEMPR7[73] ), .Y(OR4_203_Y));
    OR4 OR4_112 (.A(\R_DATA_TEMPR12[29] ), .B(\R_DATA_TEMPR13[29] ), 
        .C(\R_DATA_TEMPR14[29] ), .D(\R_DATA_TEMPR15[29] ), .Y(
        OR4_112_Y));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%12%0%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C0 (.A_DOUT({
        \R_DATA_TEMPR12[39] , \R_DATA_TEMPR12[38] , 
        \R_DATA_TEMPR12[37] , \R_DATA_TEMPR12[36] , 
        \R_DATA_TEMPR12[35] , \R_DATA_TEMPR12[34] , 
        \R_DATA_TEMPR12[33] , \R_DATA_TEMPR12[32] , 
        \R_DATA_TEMPR12[31] , \R_DATA_TEMPR12[30] , 
        \R_DATA_TEMPR12[29] , \R_DATA_TEMPR12[28] , 
        \R_DATA_TEMPR12[27] , \R_DATA_TEMPR12[26] , 
        \R_DATA_TEMPR12[25] , \R_DATA_TEMPR12[24] , 
        \R_DATA_TEMPR12[23] , \R_DATA_TEMPR12[22] , 
        \R_DATA_TEMPR12[21] , \R_DATA_TEMPR12[20] }), .B_DOUT({
        \R_DATA_TEMPR12[19] , \R_DATA_TEMPR12[18] , 
        \R_DATA_TEMPR12[17] , \R_DATA_TEMPR12[16] , 
        \R_DATA_TEMPR12[15] , \R_DATA_TEMPR12[14] , 
        \R_DATA_TEMPR12[13] , \R_DATA_TEMPR12[12] , 
        \R_DATA_TEMPR12[11] , \R_DATA_TEMPR12[10] , 
        \R_DATA_TEMPR12[9] , \R_DATA_TEMPR12[8] , \R_DATA_TEMPR12[7] , 
        \R_DATA_TEMPR12[6] , \R_DATA_TEMPR12[5] , \R_DATA_TEMPR12[4] , 
        \R_DATA_TEMPR12[3] , \R_DATA_TEMPR12[2] , \R_DATA_TEMPR12[1] , 
        \R_DATA_TEMPR12[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[12][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[3] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_204 (.A(\R_DATA_TEMPR12[8] ), .B(\R_DATA_TEMPR13[8] ), .C(
        \R_DATA_TEMPR14[8] ), .D(\R_DATA_TEMPR15[8] ), .Y(OR4_204_Y));
    OR4 OR4_84 (.A(\R_DATA_TEMPR12[34] ), .B(\R_DATA_TEMPR13[34] ), .C(
        \R_DATA_TEMPR14[34] ), .D(\R_DATA_TEMPR15[34] ), .Y(OR4_84_Y));
    OR4 OR4_42 (.A(\R_DATA_TEMPR0[52] ), .B(\R_DATA_TEMPR1[52] ), .C(
        \R_DATA_TEMPR2[52] ), .D(\R_DATA_TEMPR3[52] ), .Y(OR4_42_Y));
    OR4 OR4_190 (.A(\R_DATA_TEMPR12[46] ), .B(\R_DATA_TEMPR13[46] ), 
        .C(\R_DATA_TEMPR14[46] ), .D(\R_DATA_TEMPR15[46] ), .Y(
        OR4_190_Y));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%10%1%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C1 (.A_DOUT({
        \R_DATA_TEMPR10[79] , \R_DATA_TEMPR10[78] , 
        \R_DATA_TEMPR10[77] , \R_DATA_TEMPR10[76] , 
        \R_DATA_TEMPR10[75] , \R_DATA_TEMPR10[74] , 
        \R_DATA_TEMPR10[73] , \R_DATA_TEMPR10[72] , 
        \R_DATA_TEMPR10[71] , \R_DATA_TEMPR10[70] , 
        \R_DATA_TEMPR10[69] , \R_DATA_TEMPR10[68] , 
        \R_DATA_TEMPR10[67] , \R_DATA_TEMPR10[66] , 
        \R_DATA_TEMPR10[65] , \R_DATA_TEMPR10[64] , 
        \R_DATA_TEMPR10[63] , \R_DATA_TEMPR10[62] , 
        \R_DATA_TEMPR10[61] , \R_DATA_TEMPR10[60] }), .B_DOUT({
        \R_DATA_TEMPR10[59] , \R_DATA_TEMPR10[58] , 
        \R_DATA_TEMPR10[57] , \R_DATA_TEMPR10[56] , 
        \R_DATA_TEMPR10[55] , \R_DATA_TEMPR10[54] , 
        \R_DATA_TEMPR10[53] , \R_DATA_TEMPR10[52] , 
        \R_DATA_TEMPR10[51] , \R_DATA_TEMPR10[50] , 
        \R_DATA_TEMPR10[49] , \R_DATA_TEMPR10[48] , 
        \R_DATA_TEMPR10[47] , \R_DATA_TEMPR10[46] , 
        \R_DATA_TEMPR10[45] , \R_DATA_TEMPR10[44] , 
        \R_DATA_TEMPR10[43] , \R_DATA_TEMPR10[42] , 
        \R_DATA_TEMPR10[41] , \R_DATA_TEMPR10[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[10][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[10], \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[2] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_300 (.A(\R_DATA_TEMPR4[59] ), .B(\R_DATA_TEMPR5[59] ), .C(
        \R_DATA_TEMPR6[59] ), .D(\R_DATA_TEMPR7[59] ), .Y(OR4_300_Y));
    OR4 OR4_267 (.A(\R_DATA_TEMPR0[10] ), .B(\R_DATA_TEMPR1[10] ), .C(
        \R_DATA_TEMPR2[10] ), .D(\R_DATA_TEMPR3[10] ), .Y(OR4_267_Y));
    OR4 OR4_107 (.A(\R_DATA_TEMPR12[11] ), .B(\R_DATA_TEMPR13[11] ), 
        .C(\R_DATA_TEMPR14[11] ), .D(\R_DATA_TEMPR15[11] ), .Y(
        OR4_107_Y));
    OR4 OR4_248 (.A(\R_DATA_TEMPR8[13] ), .B(\R_DATA_TEMPR9[13] ), .C(
        \R_DATA_TEMPR10[13] ), .D(\R_DATA_TEMPR11[13] ), .Y(OR4_248_Y));
    OR4 OR4_188 (.A(\R_DATA_TEMPR8[41] ), .B(\R_DATA_TEMPR9[41] ), .C(
        \R_DATA_TEMPR10[41] ), .D(\R_DATA_TEMPR11[41] ), .Y(OR4_188_Y));
    OR4 OR4_153 (.A(\R_DATA_TEMPR12[76] ), .B(\R_DATA_TEMPR13[76] ), 
        .C(\R_DATA_TEMPR14[76] ), .D(\R_DATA_TEMPR15[76] ), .Y(
        OR4_153_Y));
    OR4 OR4_47 (.A(\R_DATA_TEMPR4[57] ), .B(\R_DATA_TEMPR5[57] ), .C(
        \R_DATA_TEMPR6[57] ), .D(\R_DATA_TEMPR7[57] ), .Y(OR4_47_Y));
    OR4 \OR4_R_DATA[6]  (.A(OR4_41_Y), .B(OR4_236_Y), .C(OR4_146_Y), 
        .D(OR4_134_Y), .Y(R_DATA[6]));
    OR4 \OR4_R_DATA[69]  (.A(OR4_56_Y), .B(OR4_15_Y), .C(OR4_249_Y), 
        .D(OR4_109_Y), .Y(R_DATA[69]));
    OR4 OR4_189 (.A(\R_DATA_TEMPR8[60] ), .B(\R_DATA_TEMPR9[60] ), .C(
        \R_DATA_TEMPR10[60] ), .D(\R_DATA_TEMPR11[60] ), .Y(OR4_189_Y));
    OR4 OR4_113 (.A(\R_DATA_TEMPR4[13] ), .B(\R_DATA_TEMPR5[13] ), .C(
        \R_DATA_TEMPR6[13] ), .D(\R_DATA_TEMPR7[13] ), .Y(OR4_113_Y));
    OR4 OR4_80 (.A(\R_DATA_TEMPR12[26] ), .B(\R_DATA_TEMPR13[26] ), .C(
        \R_DATA_TEMPR14[26] ), .D(\R_DATA_TEMPR15[26] ), .Y(OR4_80_Y));
    OR4 \OR4_R_DATA[38]  (.A(OR4_279_Y), .B(OR4_38_Y), .C(OR4_259_Y), 
        .D(OR4_171_Y), .Y(R_DATA[38]));
    OR4 \OR4_R_DATA[36]  (.A(OR4_105_Y), .B(OR4_176_Y), .C(OR4_130_Y), 
        .D(OR4_152_Y), .Y(R_DATA[36]));
    OR4 OR4_74 (.A(\R_DATA_TEMPR8[8] ), .B(\R_DATA_TEMPR9[8] ), .C(
        \R_DATA_TEMPR10[8] ), .D(\R_DATA_TEMPR11[8] ), .Y(OR4_74_Y));
    OR4 OR4_185 (.A(\R_DATA_TEMPR12[31] ), .B(\R_DATA_TEMPR13[31] ), 
        .C(\R_DATA_TEMPR14[31] ), .D(\R_DATA_TEMPR15[31] ), .Y(
        OR4_185_Y));
    OR4 \OR4_R_DATA[18]  (.A(OR4_211_Y), .B(OR4_287_Y), .C(OR4_180_Y), 
        .D(OR4_94_Y), .Y(R_DATA[18]));
    OR4 \OR4_R_DATA[16]  (.A(OR4_20_Y), .B(OR4_98_Y), .C(OR4_50_Y), .D(
        OR4_79_Y), .Y(R_DATA[16]));
    OR4 OR4_313 (.A(\R_DATA_TEMPR0[48] ), .B(\R_DATA_TEMPR1[48] ), .C(
        \R_DATA_TEMPR2[48] ), .D(\R_DATA_TEMPR3[48] ), .Y(OR4_313_Y));
    OR4 OR4_236 (.A(\R_DATA_TEMPR4[6] ), .B(\R_DATA_TEMPR5[6] ), .C(
        \R_DATA_TEMPR6[6] ), .D(\R_DATA_TEMPR7[6] ), .Y(OR4_236_Y));
    OR4 OR4_134 (.A(\R_DATA_TEMPR12[6] ), .B(\R_DATA_TEMPR13[6] ), .C(
        \R_DATA_TEMPR14[6] ), .D(\R_DATA_TEMPR15[6] ), .Y(OR4_134_Y));
    OR4 OR4_18 (.A(\R_DATA_TEMPR4[19] ), .B(\R_DATA_TEMPR5[19] ), .C(
        \R_DATA_TEMPR6[19] ), .D(\R_DATA_TEMPR7[19] ), .Y(OR4_18_Y));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%11%1%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C1 (.A_DOUT({
        \R_DATA_TEMPR11[79] , \R_DATA_TEMPR11[78] , 
        \R_DATA_TEMPR11[77] , \R_DATA_TEMPR11[76] , 
        \R_DATA_TEMPR11[75] , \R_DATA_TEMPR11[74] , 
        \R_DATA_TEMPR11[73] , \R_DATA_TEMPR11[72] , 
        \R_DATA_TEMPR11[71] , \R_DATA_TEMPR11[70] , 
        \R_DATA_TEMPR11[69] , \R_DATA_TEMPR11[68] , 
        \R_DATA_TEMPR11[67] , \R_DATA_TEMPR11[66] , 
        \R_DATA_TEMPR11[65] , \R_DATA_TEMPR11[64] , 
        \R_DATA_TEMPR11[63] , \R_DATA_TEMPR11[62] , 
        \R_DATA_TEMPR11[61] , \R_DATA_TEMPR11[60] }), .B_DOUT({
        \R_DATA_TEMPR11[59] , \R_DATA_TEMPR11[58] , 
        \R_DATA_TEMPR11[57] , \R_DATA_TEMPR11[56] , 
        \R_DATA_TEMPR11[55] , \R_DATA_TEMPR11[54] , 
        \R_DATA_TEMPR11[53] , \R_DATA_TEMPR11[52] , 
        \R_DATA_TEMPR11[51] , \R_DATA_TEMPR11[50] , 
        \R_DATA_TEMPR11[49] , \R_DATA_TEMPR11[48] , 
        \R_DATA_TEMPR11[47] , \R_DATA_TEMPR11[46] , 
        \R_DATA_TEMPR11[45] , \R_DATA_TEMPR11[44] , 
        \R_DATA_TEMPR11[43] , \R_DATA_TEMPR11[42] , 
        \R_DATA_TEMPR11[41] , \R_DATA_TEMPR11[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[11][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[2] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_68 (.A(\R_DATA_TEMPR4[34] ), .B(\R_DATA_TEMPR5[34] ), .C(
        \R_DATA_TEMPR6[34] ), .D(\R_DATA_TEMPR7[34] ), .Y(OR4_68_Y));
    OR4 OR4_208 (.A(\R_DATA_TEMPR12[57] ), .B(\R_DATA_TEMPR13[57] ), 
        .C(\R_DATA_TEMPR14[57] ), .D(\R_DATA_TEMPR15[57] ), .Y(
        OR4_208_Y));
    OR4 OR4_233 (.A(\R_DATA_TEMPR12[12] ), .B(\R_DATA_TEMPR13[12] ), 
        .C(\R_DATA_TEMPR14[12] ), .D(\R_DATA_TEMPR15[12] ), .Y(
        OR4_233_Y));
    OR4 OR4_196 (.A(\R_DATA_TEMPR8[10] ), .B(\R_DATA_TEMPR9[10] ), .C(
        \R_DATA_TEMPR10[10] ), .D(\R_DATA_TEMPR11[10] ), .Y(OR4_196_Y));
    OR4 OR4_289 (.A(\R_DATA_TEMPR12[3] ), .B(\R_DATA_TEMPR13[3] ), .C(
        \R_DATA_TEMPR14[3] ), .D(\R_DATA_TEMPR15[3] ), .Y(OR4_289_Y));
    OR4 OR4_161 (.A(\R_DATA_TEMPR12[25] ), .B(\R_DATA_TEMPR13[25] ), 
        .C(\R_DATA_TEMPR14[25] ), .D(\R_DATA_TEMPR15[25] ), .Y(
        OR4_161_Y));
    OR4 \OR4_R_DATA[41]  (.A(OR4_314_Y), .B(OR4_288_Y), .C(OR4_188_Y), 
        .D(OR4_222_Y), .Y(R_DATA[41]));
    OR4 OR4_234 (.A(\R_DATA_TEMPR12[22] ), .B(\R_DATA_TEMPR13[22] ), 
        .C(\R_DATA_TEMPR14[22] ), .D(\R_DATA_TEMPR15[22] ), .Y(
        OR4_234_Y));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%8%1%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C1 (.A_DOUT({
        \R_DATA_TEMPR8[79] , \R_DATA_TEMPR8[78] , \R_DATA_TEMPR8[77] , 
        \R_DATA_TEMPR8[76] , \R_DATA_TEMPR8[75] , \R_DATA_TEMPR8[74] , 
        \R_DATA_TEMPR8[73] , \R_DATA_TEMPR8[72] , \R_DATA_TEMPR8[71] , 
        \R_DATA_TEMPR8[70] , \R_DATA_TEMPR8[69] , \R_DATA_TEMPR8[68] , 
        \R_DATA_TEMPR8[67] , \R_DATA_TEMPR8[66] , \R_DATA_TEMPR8[65] , 
        \R_DATA_TEMPR8[64] , \R_DATA_TEMPR8[63] , \R_DATA_TEMPR8[62] , 
        \R_DATA_TEMPR8[61] , \R_DATA_TEMPR8[60] }), .B_DOUT({
        \R_DATA_TEMPR8[59] , \R_DATA_TEMPR8[58] , \R_DATA_TEMPR8[57] , 
        \R_DATA_TEMPR8[56] , \R_DATA_TEMPR8[55] , \R_DATA_TEMPR8[54] , 
        \R_DATA_TEMPR8[53] , \R_DATA_TEMPR8[52] , \R_DATA_TEMPR8[51] , 
        \R_DATA_TEMPR8[50] , \R_DATA_TEMPR8[49] , \R_DATA_TEMPR8[48] , 
        \R_DATA_TEMPR8[47] , \R_DATA_TEMPR8[46] , \R_DATA_TEMPR8[45] , 
        \R_DATA_TEMPR8[44] , \R_DATA_TEMPR8[43] , \R_DATA_TEMPR8[42] , 
        \R_DATA_TEMPR8[41] , \R_DATA_TEMPR8[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[8][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[2] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_39 (.A(\R_DATA_TEMPR4[78] ), .B(\R_DATA_TEMPR5[78] ), .C(
        \R_DATA_TEMPR6[78] ), .D(\R_DATA_TEMPR7[78] ), .Y(OR4_39_Y));
    OR4 OR4_70 (.A(\R_DATA_TEMPR8[61] ), .B(\R_DATA_TEMPR9[61] ), .C(
        \R_DATA_TEMPR10[61] ), .D(\R_DATA_TEMPR11[61] ), .Y(OR4_70_Y));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%6%0%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C0 (.A_DOUT({
        \R_DATA_TEMPR6[39] , \R_DATA_TEMPR6[38] , \R_DATA_TEMPR6[37] , 
        \R_DATA_TEMPR6[36] , \R_DATA_TEMPR6[35] , \R_DATA_TEMPR6[34] , 
        \R_DATA_TEMPR6[33] , \R_DATA_TEMPR6[32] , \R_DATA_TEMPR6[31] , 
        \R_DATA_TEMPR6[30] , \R_DATA_TEMPR6[29] , \R_DATA_TEMPR6[28] , 
        \R_DATA_TEMPR6[27] , \R_DATA_TEMPR6[26] , \R_DATA_TEMPR6[25] , 
        \R_DATA_TEMPR6[24] , \R_DATA_TEMPR6[23] , \R_DATA_TEMPR6[22] , 
        \R_DATA_TEMPR6[21] , \R_DATA_TEMPR6[20] }), .B_DOUT({
        \R_DATA_TEMPR6[19] , \R_DATA_TEMPR6[18] , \R_DATA_TEMPR6[17] , 
        \R_DATA_TEMPR6[16] , \R_DATA_TEMPR6[15] , \R_DATA_TEMPR6[14] , 
        \R_DATA_TEMPR6[13] , \R_DATA_TEMPR6[12] , \R_DATA_TEMPR6[11] , 
        \R_DATA_TEMPR6[10] , \R_DATA_TEMPR6[9] , \R_DATA_TEMPR6[8] , 
        \R_DATA_TEMPR6[7] , \R_DATA_TEMPR6[6] , \R_DATA_TEMPR6[5] , 
        \R_DATA_TEMPR6[4] , \R_DATA_TEMPR6[3] , \R_DATA_TEMPR6[2] , 
        \R_DATA_TEMPR6[1] , \R_DATA_TEMPR6[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[6][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[10], \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[1] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_306 (.A(\R_DATA_TEMPR8[34] ), .B(\R_DATA_TEMPR9[34] ), .C(
        \R_DATA_TEMPR10[34] ), .D(\R_DATA_TEMPR11[34] ), .Y(OR4_306_Y));
    OR4 OR4_308 (.A(\R_DATA_TEMPR8[45] ), .B(\R_DATA_TEMPR9[45] ), .C(
        \R_DATA_TEMPR10[45] ), .D(\R_DATA_TEMPR11[45] ), .Y(OR4_308_Y));
    OR4 OR4_137 (.A(\R_DATA_TEMPR0[75] ), .B(\R_DATA_TEMPR1[75] ), .C(
        \R_DATA_TEMPR2[75] ), .D(\R_DATA_TEMPR3[75] ), .Y(OR4_137_Y));
    OR4 OR4_251 (.A(\R_DATA_TEMPR8[57] ), .B(\R_DATA_TEMPR9[57] ), .C(
        \R_DATA_TEMPR10[57] ), .D(\R_DATA_TEMPR11[57] ), .Y(OR4_251_Y));
    OR4 \OR4_R_DATA[5]  (.A(OR4_114_Y), .B(OR4_256_Y), .C(OR4_175_Y), 
        .D(OR4_10_Y), .Y(R_DATA[5]));
    OR4 OR4_227 (.A(\R_DATA_TEMPR8[14] ), .B(\R_DATA_TEMPR9[14] ), .C(
        \R_DATA_TEMPR10[14] ), .D(\R_DATA_TEMPR11[14] ), .Y(OR4_227_Y));
    OR4 OR4_140 (.A(\R_DATA_TEMPR0[46] ), .B(\R_DATA_TEMPR1[46] ), .C(
        \R_DATA_TEMPR2[46] ), .D(\R_DATA_TEMPR3[46] ), .Y(OR4_140_Y));
    OR4 OR4_55 (.A(\R_DATA_TEMPR0[65] ), .B(\R_DATA_TEMPR1[65] ), .C(
        \R_DATA_TEMPR2[65] ), .D(\R_DATA_TEMPR3[65] ), .Y(OR4_55_Y));
    OR4 \OR4_R_DATA[79]  (.A(OR4_139_Y), .B(OR4_103_Y), .C(OR4_9_Y), 
        .D(OR4_197_Y), .Y(R_DATA[79]));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%15%0%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C0 (.A_DOUT({
        \R_DATA_TEMPR15[39] , \R_DATA_TEMPR15[38] , 
        \R_DATA_TEMPR15[37] , \R_DATA_TEMPR15[36] , 
        \R_DATA_TEMPR15[35] , \R_DATA_TEMPR15[34] , 
        \R_DATA_TEMPR15[33] , \R_DATA_TEMPR15[32] , 
        \R_DATA_TEMPR15[31] , \R_DATA_TEMPR15[30] , 
        \R_DATA_TEMPR15[29] , \R_DATA_TEMPR15[28] , 
        \R_DATA_TEMPR15[27] , \R_DATA_TEMPR15[26] , 
        \R_DATA_TEMPR15[25] , \R_DATA_TEMPR15[24] , 
        \R_DATA_TEMPR15[23] , \R_DATA_TEMPR15[22] , 
        \R_DATA_TEMPR15[21] , \R_DATA_TEMPR15[20] }), .B_DOUT({
        \R_DATA_TEMPR15[19] , \R_DATA_TEMPR15[18] , 
        \R_DATA_TEMPR15[17] , \R_DATA_TEMPR15[16] , 
        \R_DATA_TEMPR15[15] , \R_DATA_TEMPR15[14] , 
        \R_DATA_TEMPR15[13] , \R_DATA_TEMPR15[12] , 
        \R_DATA_TEMPR15[11] , \R_DATA_TEMPR15[10] , 
        \R_DATA_TEMPR15[9] , \R_DATA_TEMPR15[8] , \R_DATA_TEMPR15[7] , 
        \R_DATA_TEMPR15[6] , \R_DATA_TEMPR15[5] , \R_DATA_TEMPR15[4] , 
        \R_DATA_TEMPR15[3] , \R_DATA_TEMPR15[2] , \R_DATA_TEMPR15[1] , 
        \R_DATA_TEMPR15[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[15][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[3] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[3] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_95 (.A(\R_DATA_TEMPR4[27] ), .B(\R_DATA_TEMPR5[27] ), .C(
        \R_DATA_TEMPR6[27] ), .D(\R_DATA_TEMPR7[27] ), .Y(OR4_95_Y));
    OR4 OR4_211 (.A(\R_DATA_TEMPR0[18] ), .B(\R_DATA_TEMPR1[18] ), .C(
        \R_DATA_TEMPR2[18] ), .D(\R_DATA_TEMPR3[18] ), .Y(OR4_211_Y));
    OR4 OR4_168 (.A(\R_DATA_TEMPR4[37] ), .B(\R_DATA_TEMPR5[37] ), .C(
        \R_DATA_TEMPR6[37] ), .D(\R_DATA_TEMPR7[37] ), .Y(OR4_168_Y));
    OR4 \OR4_R_DATA[67]  (.A(OR4_276_Y), .B(OR4_88_Y), .C(OR4_291_Y), 
        .D(OR4_237_Y), .Y(R_DATA[67]));
    OR4 OR4_277 (.A(\R_DATA_TEMPR0[13] ), .B(\R_DATA_TEMPR1[13] ), .C(
        \R_DATA_TEMPR2[13] ), .D(\R_DATA_TEMPR3[13] ), .Y(OR4_277_Y));
    OR4 OR4_51 (.A(\R_DATA_TEMPR8[37] ), .B(\R_DATA_TEMPR9[37] ), .C(
        \R_DATA_TEMPR10[37] ), .D(\R_DATA_TEMPR11[37] ), .Y(OR4_51_Y));
    OR4 OR4_83 (.A(\R_DATA_TEMPR8[52] ), .B(\R_DATA_TEMPR9[52] ), .C(
        \R_DATA_TEMPR10[52] ), .D(\R_DATA_TEMPR11[52] ), .Y(OR4_83_Y));
    OR4 OR4_91 (.A(\R_DATA_TEMPR4[42] ), .B(\R_DATA_TEMPR5[42] ), .C(
        \R_DATA_TEMPR6[42] ), .D(\R_DATA_TEMPR7[42] ), .Y(OR4_91_Y));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%4%1%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C1 (.A_DOUT({
        \R_DATA_TEMPR4[79] , \R_DATA_TEMPR4[78] , \R_DATA_TEMPR4[77] , 
        \R_DATA_TEMPR4[76] , \R_DATA_TEMPR4[75] , \R_DATA_TEMPR4[74] , 
        \R_DATA_TEMPR4[73] , \R_DATA_TEMPR4[72] , \R_DATA_TEMPR4[71] , 
        \R_DATA_TEMPR4[70] , \R_DATA_TEMPR4[69] , \R_DATA_TEMPR4[68] , 
        \R_DATA_TEMPR4[67] , \R_DATA_TEMPR4[66] , \R_DATA_TEMPR4[65] , 
        \R_DATA_TEMPR4[64] , \R_DATA_TEMPR4[63] , \R_DATA_TEMPR4[62] , 
        \R_DATA_TEMPR4[61] , \R_DATA_TEMPR4[60] }), .B_DOUT({
        \R_DATA_TEMPR4[59] , \R_DATA_TEMPR4[58] , \R_DATA_TEMPR4[57] , 
        \R_DATA_TEMPR4[56] , \R_DATA_TEMPR4[55] , \R_DATA_TEMPR4[54] , 
        \R_DATA_TEMPR4[53] , \R_DATA_TEMPR4[52] , \R_DATA_TEMPR4[51] , 
        \R_DATA_TEMPR4[50] , \R_DATA_TEMPR4[49] , \R_DATA_TEMPR4[48] , 
        \R_DATA_TEMPR4[47] , \R_DATA_TEMPR4[46] , \R_DATA_TEMPR4[45] , 
        \R_DATA_TEMPR4[44] , \R_DATA_TEMPR4[43] , \R_DATA_TEMPR4[42] , 
        \R_DATA_TEMPR4[41] , \R_DATA_TEMPR4[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[4][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[1] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[9]  (.A(OR4_46_Y), .B(OR4_305_Y), .C(OR4_221_Y), 
        .D(OR4_218_Y), .Y(R_DATA[9]));
    OR4 OR4_169 (.A(\R_DATA_TEMPR4[77] ), .B(\R_DATA_TEMPR5[77] ), .C(
        \R_DATA_TEMPR6[77] ), .D(\R_DATA_TEMPR7[77] ), .Y(OR4_169_Y));
    OR4 \OR4_R_DATA[58]  (.A(OR4_155_Y), .B(OR4_240_Y), .C(OR4_141_Y), 
        .D(OR4_48_Y), .Y(R_DATA[58]));
    OR4 \OR4_R_DATA[56]  (.A(OR4_302_Y), .B(OR4_58_Y), .C(OR4_7_Y), .D(
        OR4_27_Y), .Y(R_DATA[56]));
    OR4 OR4_8 (.A(\R_DATA_TEMPR8[39] ), .B(\R_DATA_TEMPR9[39] ), .C(
        \R_DATA_TEMPR10[39] ), .D(\R_DATA_TEMPR11[39] ), .Y(OR4_8_Y));
    OR4 OR4_100 (.A(\R_DATA_TEMPR4[26] ), .B(\R_DATA_TEMPR5[26] ), .C(
        \R_DATA_TEMPR6[26] ), .D(\R_DATA_TEMPR7[26] ), .Y(OR4_100_Y));
    OR4 OR4_238 (.A(\R_DATA_TEMPR0[57] ), .B(\R_DATA_TEMPR1[57] ), .C(
        \R_DATA_TEMPR2[57] ), .D(\R_DATA_TEMPR3[57] ), .Y(OR4_238_Y));
    OR4 \OR4_R_DATA[44]  (.A(OR4_301_Y), .B(OR4_101_Y), .C(OR4_16_Y), 
        .D(OR4_119_Y), .Y(R_DATA[44]));
    OR4 OR4_295 (.A(\R_DATA_TEMPR12[43] ), .B(\R_DATA_TEMPR13[43] ), 
        .C(\R_DATA_TEMPR14[43] ), .D(\R_DATA_TEMPR15[43] ), .Y(
        OR4_295_Y));
    OR4 OR4_286 (.A(\R_DATA_TEMPR0[71] ), .B(\R_DATA_TEMPR1[71] ), .C(
        \R_DATA_TEMPR2[71] ), .D(\R_DATA_TEMPR3[71] ), .Y(OR4_286_Y));
    OR4 OR4_165 (.A(\R_DATA_TEMPR0[72] ), .B(\R_DATA_TEMPR1[72] ), .C(
        \R_DATA_TEMPR2[72] ), .D(\R_DATA_TEMPR3[72] ), .Y(OR4_165_Y));
    OR4 OR4_29 (.A(\R_DATA_TEMPR12[60] ), .B(\R_DATA_TEMPR13[60] ), .C(
        \R_DATA_TEMPR14[60] ), .D(\R_DATA_TEMPR15[60] ), .Y(OR4_29_Y));
    OR4 \OR4_R_DATA[43]  (.A(OR4_77_Y), .B(OR4_229_Y), .C(OR4_32_Y), 
        .D(OR4_295_Y), .Y(R_DATA[43]));
    OR4 OR4_184 (.A(\R_DATA_TEMPR8[54] ), .B(\R_DATA_TEMPR9[54] ), .C(
        \R_DATA_TEMPR10[54] ), .D(\R_DATA_TEMPR11[54] ), .Y(OR4_184_Y));
    OR4 OR4_283 (.A(\R_DATA_TEMPR12[54] ), .B(\R_DATA_TEMPR13[54] ), 
        .C(\R_DATA_TEMPR14[54] ), .D(\R_DATA_TEMPR15[54] ), .Y(
        OR4_283_Y));
    OR4 OR4_146 (.A(\R_DATA_TEMPR8[6] ), .B(\R_DATA_TEMPR9[6] ), .C(
        \R_DATA_TEMPR10[6] ), .D(\R_DATA_TEMPR11[6] ), .Y(OR4_146_Y));
    OR4 OR4_66 (.A(\R_DATA_TEMPR0[40] ), .B(\R_DATA_TEMPR1[40] ), .C(
        \R_DATA_TEMPR2[40] ), .D(\R_DATA_TEMPR3[40] ), .Y(OR4_66_Y));
    OR4 OR4_16 (.A(\R_DATA_TEMPR8[44] ), .B(\R_DATA_TEMPR9[44] ), .C(
        \R_DATA_TEMPR10[44] ), .D(\R_DATA_TEMPR11[44] ), .Y(OR4_16_Y));
    OR4 OR4_121 (.A(\R_DATA_TEMPR12[70] ), .B(\R_DATA_TEMPR13[70] ), 
        .C(\R_DATA_TEMPR14[70] ), .D(\R_DATA_TEMPR15[70] ), .Y(
        OR4_121_Y));
    OR4 OR4_45 (.A(\R_DATA_TEMPR4[25] ), .B(\R_DATA_TEMPR5[25] ), .C(
        \R_DATA_TEMPR6[25] ), .D(\R_DATA_TEMPR7[25] ), .Y(OR4_45_Y));
    OR4 \OR4_R_DATA[60]  (.A(OR4_263_Y), .B(OR4_49_Y), .C(OR4_189_Y), 
        .D(OR4_29_Y), .Y(R_DATA[60]));
    OR4 OR4_73 (.A(\R_DATA_TEMPR8[11] ), .B(\R_DATA_TEMPR9[11] ), .C(
        \R_DATA_TEMPR10[11] ), .D(\R_DATA_TEMPR11[11] ), .Y(OR4_73_Y));
    OR4 OR4_284 (.A(\R_DATA_TEMPR0[31] ), .B(\R_DATA_TEMPR1[31] ), .C(
        \R_DATA_TEMPR2[31] ), .D(\R_DATA_TEMPR3[31] ), .Y(OR4_284_Y));
    OR4 OR4_269 (.A(\R_DATA_TEMPR8[30] ), .B(\R_DATA_TEMPR9[30] ), .C(
        \R_DATA_TEMPR10[30] ), .D(\R_DATA_TEMPR11[30] ), .Y(OR4_269_Y));
    OR4 \OR4_R_DATA[45]  (.A(OR4_167_Y), .B(OR4_156_Y), .C(OR4_308_Y), 
        .D(OR4_275_Y), .Y(R_DATA[45]));
    OR4 OR4_34 (.A(\R_DATA_TEMPR12[10] ), .B(\R_DATA_TEMPR13[10] ), .C(
        \R_DATA_TEMPR14[10] ), .D(\R_DATA_TEMPR15[10] ), .Y(OR4_34_Y));
    OR4 OR4_290 (.A(\R_DATA_TEMPR4[28] ), .B(\R_DATA_TEMPR5[28] ), .C(
        \R_DATA_TEMPR6[28] ), .D(\R_DATA_TEMPR7[28] ), .Y(OR4_290_Y));
    OR4 OR4_171 (.A(\R_DATA_TEMPR12[38] ), .B(\R_DATA_TEMPR13[38] ), 
        .C(\R_DATA_TEMPR14[38] ), .D(\R_DATA_TEMPR15[38] ), .Y(
        OR4_171_Y));
    OR4 OR4_41 (.A(\R_DATA_TEMPR0[6] ), .B(\R_DATA_TEMPR1[6] ), .C(
        \R_DATA_TEMPR2[6] ), .D(\R_DATA_TEMPR3[6] ), .Y(OR4_41_Y));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%1%1%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C1 (.A_DOUT({
        \R_DATA_TEMPR1[79] , \R_DATA_TEMPR1[78] , \R_DATA_TEMPR1[77] , 
        \R_DATA_TEMPR1[76] , \R_DATA_TEMPR1[75] , \R_DATA_TEMPR1[74] , 
        \R_DATA_TEMPR1[73] , \R_DATA_TEMPR1[72] , \R_DATA_TEMPR1[71] , 
        \R_DATA_TEMPR1[70] , \R_DATA_TEMPR1[69] , \R_DATA_TEMPR1[68] , 
        \R_DATA_TEMPR1[67] , \R_DATA_TEMPR1[66] , \R_DATA_TEMPR1[65] , 
        \R_DATA_TEMPR1[64] , \R_DATA_TEMPR1[63] , \R_DATA_TEMPR1[62] , 
        \R_DATA_TEMPR1[61] , \R_DATA_TEMPR1[60] }), .B_DOUT({
        \R_DATA_TEMPR1[59] , \R_DATA_TEMPR1[58] , \R_DATA_TEMPR1[57] , 
        \R_DATA_TEMPR1[56] , \R_DATA_TEMPR1[55] , \R_DATA_TEMPR1[54] , 
        \R_DATA_TEMPR1[53] , \R_DATA_TEMPR1[52] , \R_DATA_TEMPR1[51] , 
        \R_DATA_TEMPR1[50] , \R_DATA_TEMPR1[49] , \R_DATA_TEMPR1[48] , 
        \R_DATA_TEMPR1[47] , \R_DATA_TEMPR1[46] , \R_DATA_TEMPR1[45] , 
        \R_DATA_TEMPR1[44] , \R_DATA_TEMPR1[43] , \R_DATA_TEMPR1[42] , 
        \R_DATA_TEMPR1[41] , \R_DATA_TEMPR1[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[1][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[0] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_7 (.A(\R_DATA_TEMPR8[56] ), .B(\R_DATA_TEMPR9[56] ), .C(
        \R_DATA_TEMPR10[56] ), .D(\R_DATA_TEMPR11[56] ), .Y(OR4_7_Y));
    OR4 OR4_187 (.A(\R_DATA_TEMPR0[64] ), .B(\R_DATA_TEMPR1[64] ), .C(
        \R_DATA_TEMPR2[64] ), .D(\R_DATA_TEMPR3[64] ), .Y(OR4_187_Y));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%0%0%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C0 (.A_DOUT({
        \R_DATA_TEMPR0[39] , \R_DATA_TEMPR0[38] , \R_DATA_TEMPR0[37] , 
        \R_DATA_TEMPR0[36] , \R_DATA_TEMPR0[35] , \R_DATA_TEMPR0[34] , 
        \R_DATA_TEMPR0[33] , \R_DATA_TEMPR0[32] , \R_DATA_TEMPR0[31] , 
        \R_DATA_TEMPR0[30] , \R_DATA_TEMPR0[29] , \R_DATA_TEMPR0[28] , 
        \R_DATA_TEMPR0[27] , \R_DATA_TEMPR0[26] , \R_DATA_TEMPR0[25] , 
        \R_DATA_TEMPR0[24] , \R_DATA_TEMPR0[23] , \R_DATA_TEMPR0[22] , 
        \R_DATA_TEMPR0[21] , \R_DATA_TEMPR0[20] }), .B_DOUT({
        \R_DATA_TEMPR0[19] , \R_DATA_TEMPR0[18] , \R_DATA_TEMPR0[17] , 
        \R_DATA_TEMPR0[16] , \R_DATA_TEMPR0[15] , \R_DATA_TEMPR0[14] , 
        \R_DATA_TEMPR0[13] , \R_DATA_TEMPR0[12] , \R_DATA_TEMPR0[11] , 
        \R_DATA_TEMPR0[10] , \R_DATA_TEMPR0[9] , \R_DATA_TEMPR0[8] , 
        \R_DATA_TEMPR0[7] , \R_DATA_TEMPR0[6] , \R_DATA_TEMPR0[5] , 
        \R_DATA_TEMPR0[4] , \R_DATA_TEMPR0[3] , \R_DATA_TEMPR0[2] , 
        \R_DATA_TEMPR0[1] , \R_DATA_TEMPR0[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[0][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[0] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%0%1%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C1 (.A_DOUT({
        \R_DATA_TEMPR0[79] , \R_DATA_TEMPR0[78] , \R_DATA_TEMPR0[77] , 
        \R_DATA_TEMPR0[76] , \R_DATA_TEMPR0[75] , \R_DATA_TEMPR0[74] , 
        \R_DATA_TEMPR0[73] , \R_DATA_TEMPR0[72] , \R_DATA_TEMPR0[71] , 
        \R_DATA_TEMPR0[70] , \R_DATA_TEMPR0[69] , \R_DATA_TEMPR0[68] , 
        \R_DATA_TEMPR0[67] , \R_DATA_TEMPR0[66] , \R_DATA_TEMPR0[65] , 
        \R_DATA_TEMPR0[64] , \R_DATA_TEMPR0[63] , \R_DATA_TEMPR0[62] , 
        \R_DATA_TEMPR0[61] , \R_DATA_TEMPR0[60] }), .B_DOUT({
        \R_DATA_TEMPR0[59] , \R_DATA_TEMPR0[58] , \R_DATA_TEMPR0[57] , 
        \R_DATA_TEMPR0[56] , \R_DATA_TEMPR0[55] , \R_DATA_TEMPR0[54] , 
        \R_DATA_TEMPR0[53] , \R_DATA_TEMPR0[52] , \R_DATA_TEMPR0[51] , 
        \R_DATA_TEMPR0[50] , \R_DATA_TEMPR0[49] , \R_DATA_TEMPR0[48] , 
        \R_DATA_TEMPR0[47] , \R_DATA_TEMPR0[46] , \R_DATA_TEMPR0[45] , 
        \R_DATA_TEMPR0[44] , \R_DATA_TEMPR0[43] , \R_DATA_TEMPR0[42] , 
        \R_DATA_TEMPR0[41] , \R_DATA_TEMPR0[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[0][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[0] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[77]  (.A(OR4_35_Y), .B(OR4_169_Y), .C(OR4_52_Y), 
        .D(OR4_318_Y), .Y(R_DATA[77]));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%3%0%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C0 (.A_DOUT({
        \R_DATA_TEMPR3[39] , \R_DATA_TEMPR3[38] , \R_DATA_TEMPR3[37] , 
        \R_DATA_TEMPR3[36] , \R_DATA_TEMPR3[35] , \R_DATA_TEMPR3[34] , 
        \R_DATA_TEMPR3[33] , \R_DATA_TEMPR3[32] , \R_DATA_TEMPR3[31] , 
        \R_DATA_TEMPR3[30] , \R_DATA_TEMPR3[29] , \R_DATA_TEMPR3[28] , 
        \R_DATA_TEMPR3[27] , \R_DATA_TEMPR3[26] , \R_DATA_TEMPR3[25] , 
        \R_DATA_TEMPR3[24] , \R_DATA_TEMPR3[23] , \R_DATA_TEMPR3[22] , 
        \R_DATA_TEMPR3[21] , \R_DATA_TEMPR3[20] }), .B_DOUT({
        \R_DATA_TEMPR3[19] , \R_DATA_TEMPR3[18] , \R_DATA_TEMPR3[17] , 
        \R_DATA_TEMPR3[16] , \R_DATA_TEMPR3[15] , \R_DATA_TEMPR3[14] , 
        \R_DATA_TEMPR3[13] , \R_DATA_TEMPR3[12] , \R_DATA_TEMPR3[11] , 
        \R_DATA_TEMPR3[10] , \R_DATA_TEMPR3[9] , \R_DATA_TEMPR3[8] , 
        \R_DATA_TEMPR3[7] , \R_DATA_TEMPR3[6] , \R_DATA_TEMPR3[5] , 
        \R_DATA_TEMPR3[4] , \R_DATA_TEMPR3[3] , \R_DATA_TEMPR3[2] , 
        \R_DATA_TEMPR3[1] , \R_DATA_TEMPR3[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[3][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[0] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_106 (.A(\R_DATA_TEMPR0[76] ), .B(\R_DATA_TEMPR1[76] ), .C(
        \R_DATA_TEMPR2[76] ), .D(\R_DATA_TEMPR3[76] ), .Y(OR4_106_Y));
    OR4 OR4_128 (.A(\R_DATA_TEMPR0[3] ), .B(\R_DATA_TEMPR1[3] ), .C(
        \R_DATA_TEMPR2[3] ), .D(\R_DATA_TEMPR3[3] ), .Y(OR4_128_Y));
    OR4 \OR4_R_DATA[42]  (.A(OR4_210_Y), .B(OR4_91_Y), .C(OR4_232_Y), 
        .D(OR4_24_Y), .Y(R_DATA[42]));
    CFG3 #( .INIT(8'h40) )  \CFG3_BLKY2[1]  (.A(R_ADDR[12]), .B(
        R_ADDR[11]), .C(R_EN), .Y(\BLKY2[1] ));
    OR4 OR4_30 (.A(\R_DATA_TEMPR0[33] ), .B(\R_DATA_TEMPR1[33] ), .C(
        \R_DATA_TEMPR2[33] ), .D(\R_DATA_TEMPR3[33] ), .Y(OR4_30_Y));
    OR4 OR4_88 (.A(\R_DATA_TEMPR4[67] ), .B(\R_DATA_TEMPR5[67] ), .C(
        \R_DATA_TEMPR6[67] ), .D(\R_DATA_TEMPR7[67] ), .Y(OR4_88_Y));
    CFG3 #( .INIT(8'h80) )  \CFG3_BLKY2[3]  (.A(R_ADDR[12]), .B(
        R_ADDR[11]), .C(R_EN), .Y(\BLKY2[3] ));
    OR4 OR4_292 (.A(\R_DATA_TEMPR8[17] ), .B(\R_DATA_TEMPR9[17] ), .C(
        \R_DATA_TEMPR10[17] ), .D(\R_DATA_TEMPR11[17] ), .Y(OR4_292_Y));
    OR4 OR4_130 (.A(\R_DATA_TEMPR8[36] ), .B(\R_DATA_TEMPR9[36] ), .C(
        \R_DATA_TEMPR10[36] ), .D(\R_DATA_TEMPR11[36] ), .Y(OR4_130_Y));
    OR4 OR4_129 (.A(\R_DATA_TEMPR4[51] ), .B(\R_DATA_TEMPR5[51] ), .C(
        \R_DATA_TEMPR6[51] ), .D(\R_DATA_TEMPR7[51] ), .Y(OR4_129_Y));
    OR4 OR4_178 (.A(\R_DATA_TEMPR8[68] ), .B(\R_DATA_TEMPR9[68] ), .C(
        \R_DATA_TEMPR10[68] ), .D(\R_DATA_TEMPR11[68] ), .Y(OR4_178_Y));
    OR4 OR4_192 (.A(\R_DATA_TEMPR0[14] ), .B(\R_DATA_TEMPR1[14] ), .C(
        \R_DATA_TEMPR2[14] ), .D(\R_DATA_TEMPR3[14] ), .Y(OR4_192_Y));
    OR4 OR4_314 (.A(\R_DATA_TEMPR0[41] ), .B(\R_DATA_TEMPR1[41] ), .C(
        \R_DATA_TEMPR2[41] ), .D(\R_DATA_TEMPR3[41] ), .Y(OR4_314_Y));
    OR4 OR4_302 (.A(\R_DATA_TEMPR0[56] ), .B(\R_DATA_TEMPR1[56] ), .C(
        \R_DATA_TEMPR2[56] ), .D(\R_DATA_TEMPR3[56] ), .Y(OR4_302_Y));
    OR4 OR4_288 (.A(\R_DATA_TEMPR4[41] ), .B(\R_DATA_TEMPR5[41] ), .C(
        \R_DATA_TEMPR6[41] ), .D(\R_DATA_TEMPR7[41] ), .Y(OR4_288_Y));
    OR4 OR4_125 (.A(\R_DATA_TEMPR4[35] ), .B(\R_DATA_TEMPR5[35] ), .C(
        \R_DATA_TEMPR6[35] ), .D(\R_DATA_TEMPR7[35] ), .Y(OR4_125_Y));
    OR4 \OR4_R_DATA[70]  (.A(OR4_23_Y), .B(OR4_133_Y), .C(OR4_271_Y), 
        .D(OR4_121_Y), .Y(R_DATA[70]));
    OR4 OR4_245 (.A(\R_DATA_TEMPR12[75] ), .B(\R_DATA_TEMPR13[75] ), 
        .C(\R_DATA_TEMPR14[75] ), .D(\R_DATA_TEMPR15[75] ), .Y(
        OR4_245_Y));
    OR4 \OR4_R_DATA[31]  (.A(OR4_284_Y), .B(OR4_252_Y), .C(OR4_149_Y), 
        .D(OR4_185_Y), .Y(R_DATA[31]));
    OR4 OR4_24 (.A(\R_DATA_TEMPR12[42] ), .B(\R_DATA_TEMPR13[42] ), .C(
        \R_DATA_TEMPR14[42] ), .D(\R_DATA_TEMPR15[42] ), .Y(OR4_24_Y));
    OR4 OR4_179 (.A(\R_DATA_TEMPR12[63] ), .B(\R_DATA_TEMPR13[63] ), 
        .C(\R_DATA_TEMPR14[63] ), .D(\R_DATA_TEMPR15[63] ), .Y(
        OR4_179_Y));
    OR4 OR4_12 (.A(\R_DATA_TEMPR12[4] ), .B(\R_DATA_TEMPR13[4] ), .C(
        \R_DATA_TEMPR14[4] ), .D(\R_DATA_TEMPR15[4] ), .Y(OR4_12_Y));
    OR4 OR4_62 (.A(\R_DATA_TEMPR0[15] ), .B(\R_DATA_TEMPR1[15] ), .C(
        \R_DATA_TEMPR2[15] ), .D(\R_DATA_TEMPR3[15] ), .Y(OR4_62_Y));
    OR4 OR4_266 (.A(\R_DATA_TEMPR0[74] ), .B(\R_DATA_TEMPR1[74] ), .C(
        \R_DATA_TEMPR2[74] ), .D(\R_DATA_TEMPR3[74] ), .Y(OR4_266_Y));
    OR4 \OR4_R_DATA[11]  (.A(OR4_215_Y), .B(OR4_173_Y), .C(OR4_73_Y), 
        .D(OR4_107_Y), .Y(R_DATA[11]));
    OR4 OR4_164 (.A(\R_DATA_TEMPR0[32] ), .B(\R_DATA_TEMPR1[32] ), .C(
        \R_DATA_TEMPR2[32] ), .D(\R_DATA_TEMPR3[32] ), .Y(OR4_164_Y));
    OR4 OR4_311 (.A(\R_DATA_TEMPR12[32] ), .B(\R_DATA_TEMPR13[32] ), 
        .C(\R_DATA_TEMPR14[32] ), .D(\R_DATA_TEMPR15[32] ), .Y(
        OR4_311_Y));
    OR4 OR4_263 (.A(\R_DATA_TEMPR0[60] ), .B(\R_DATA_TEMPR1[60] ), .C(
        \R_DATA_TEMPR2[60] ), .D(\R_DATA_TEMPR3[60] ), .Y(OR4_263_Y));
    OR4 OR4_257 (.A(\R_DATA_TEMPR4[52] ), .B(\R_DATA_TEMPR5[52] ), .C(
        \R_DATA_TEMPR6[52] ), .D(\R_DATA_TEMPR7[52] ), .Y(OR4_257_Y));
    OR4 OR4_229 (.A(\R_DATA_TEMPR4[43] ), .B(\R_DATA_TEMPR5[43] ), .C(
        \R_DATA_TEMPR6[43] ), .D(\R_DATA_TEMPR7[43] ), .Y(OR4_229_Y));
    OR4 OR4_175 (.A(\R_DATA_TEMPR8[5] ), .B(\R_DATA_TEMPR9[5] ), .C(
        \R_DATA_TEMPR10[5] ), .D(\R_DATA_TEMPR11[5] ), .Y(OR4_175_Y));
    OR4 \OR4_R_DATA[29]  (.A(OR4_65_Y), .B(OR4_19_Y), .C(OR4_255_Y), 
        .D(OR4_112_Y), .Y(R_DATA[29]));
    OR4 OR4_78 (.A(\R_DATA_TEMPR8[21] ), .B(\R_DATA_TEMPR9[21] ), .C(
        \R_DATA_TEMPR10[21] ), .D(\R_DATA_TEMPR11[21] ), .Y(OR4_78_Y));
    OR4 OR4_67 (.A(\R_DATA_TEMPR12[51] ), .B(\R_DATA_TEMPR13[51] ), .C(
        \R_DATA_TEMPR14[51] ), .D(\R_DATA_TEMPR15[51] ), .Y(OR4_67_Y));
    OR4 OR4_17 (.A(\R_DATA_TEMPR0[66] ), .B(\R_DATA_TEMPR1[66] ), .C(
        \R_DATA_TEMPR2[66] ), .D(\R_DATA_TEMPR3[66] ), .Y(OR4_17_Y));
    OR4 OR4_264 (.A(\R_DATA_TEMPR4[54] ), .B(\R_DATA_TEMPR5[54] ), .C(
        \R_DATA_TEMPR6[54] ), .D(\R_DATA_TEMPR7[54] ), .Y(OR4_264_Y));
    OR4 OR4_240 (.A(\R_DATA_TEMPR4[58] ), .B(\R_DATA_TEMPR5[58] ), .C(
        \R_DATA_TEMPR6[58] ), .D(\R_DATA_TEMPR7[58] ), .Y(OR4_240_Y));
    OR4 OR4_217 (.A(\R_DATA_TEMPR0[21] ), .B(\R_DATA_TEMPR1[21] ), .C(
        \R_DATA_TEMPR2[21] ), .D(\R_DATA_TEMPR3[21] ), .Y(OR4_217_Y));
    OR4 OR4_279 (.A(\R_DATA_TEMPR0[38] ), .B(\R_DATA_TEMPR1[38] ), .C(
        \R_DATA_TEMPR2[38] ), .D(\R_DATA_TEMPR3[38] ), .Y(OR4_279_Y));
    OR4 OR4_136 (.A(\R_DATA_TEMPR0[35] ), .B(\R_DATA_TEMPR1[35] ), .C(
        \R_DATA_TEMPR2[35] ), .D(\R_DATA_TEMPR3[35] ), .Y(OR4_136_Y));
    OR4 OR4_205 (.A(\R_DATA_TEMPR0[68] ), .B(\R_DATA_TEMPR1[68] ), .C(
        \R_DATA_TEMPR2[68] ), .D(\R_DATA_TEMPR3[68] ), .Y(OR4_205_Y));
    OR4 OR4_20 (.A(\R_DATA_TEMPR0[16] ), .B(\R_DATA_TEMPR1[16] ), .C(
        \R_DATA_TEMPR2[16] ), .D(\R_DATA_TEMPR3[16] ), .Y(OR4_20_Y));
    OR4 OR4_193 (.A(\R_DATA_TEMPR8[65] ), .B(\R_DATA_TEMPR9[65] ), .C(
        \R_DATA_TEMPR10[65] ), .D(\R_DATA_TEMPR11[65] ), .Y(OR4_193_Y));
    OR4 OR4_167 (.A(\R_DATA_TEMPR0[45] ), .B(\R_DATA_TEMPR1[45] ), .C(
        \R_DATA_TEMPR2[45] ), .D(\R_DATA_TEMPR3[45] ), .Y(OR4_167_Y));
    OR4 OR4_33 (.A(\R_DATA_TEMPR0[37] ), .B(\R_DATA_TEMPR1[37] ), .C(
        \R_DATA_TEMPR2[37] ), .D(\R_DATA_TEMPR3[37] ), .Y(OR4_33_Y));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%12%1%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C1 (.A_DOUT({
        \R_DATA_TEMPR12[79] , \R_DATA_TEMPR12[78] , 
        \R_DATA_TEMPR12[77] , \R_DATA_TEMPR12[76] , 
        \R_DATA_TEMPR12[75] , \R_DATA_TEMPR12[74] , 
        \R_DATA_TEMPR12[73] , \R_DATA_TEMPR12[72] , 
        \R_DATA_TEMPR12[71] , \R_DATA_TEMPR12[70] , 
        \R_DATA_TEMPR12[69] , \R_DATA_TEMPR12[68] , 
        \R_DATA_TEMPR12[67] , \R_DATA_TEMPR12[66] , 
        \R_DATA_TEMPR12[65] , \R_DATA_TEMPR12[64] , 
        \R_DATA_TEMPR12[63] , \R_DATA_TEMPR12[62] , 
        \R_DATA_TEMPR12[61] , \R_DATA_TEMPR12[60] }), .B_DOUT({
        \R_DATA_TEMPR12[59] , \R_DATA_TEMPR12[58] , 
        \R_DATA_TEMPR12[57] , \R_DATA_TEMPR12[56] , 
        \R_DATA_TEMPR12[55] , \R_DATA_TEMPR12[54] , 
        \R_DATA_TEMPR12[53] , \R_DATA_TEMPR12[52] , 
        \R_DATA_TEMPR12[51] , \R_DATA_TEMPR12[50] , 
        \R_DATA_TEMPR12[49] , \R_DATA_TEMPR12[48] , 
        \R_DATA_TEMPR12[47] , \R_DATA_TEMPR12[46] , 
        \R_DATA_TEMPR12[45] , \R_DATA_TEMPR12[44] , 
        \R_DATA_TEMPR12[43] , \R_DATA_TEMPR12[42] , 
        \R_DATA_TEMPR12[41] , \R_DATA_TEMPR12[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[12][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[3] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%11%0%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C0 (.A_DOUT({
        \R_DATA_TEMPR11[39] , \R_DATA_TEMPR11[38] , 
        \R_DATA_TEMPR11[37] , \R_DATA_TEMPR11[36] , 
        \R_DATA_TEMPR11[35] , \R_DATA_TEMPR11[34] , 
        \R_DATA_TEMPR11[33] , \R_DATA_TEMPR11[32] , 
        \R_DATA_TEMPR11[31] , \R_DATA_TEMPR11[30] , 
        \R_DATA_TEMPR11[29] , \R_DATA_TEMPR11[28] , 
        \R_DATA_TEMPR11[27] , \R_DATA_TEMPR11[26] , 
        \R_DATA_TEMPR11[25] , \R_DATA_TEMPR11[24] , 
        \R_DATA_TEMPR11[23] , \R_DATA_TEMPR11[22] , 
        \R_DATA_TEMPR11[21] , \R_DATA_TEMPR11[20] }), .B_DOUT({
        \R_DATA_TEMPR11[19] , \R_DATA_TEMPR11[18] , 
        \R_DATA_TEMPR11[17] , \R_DATA_TEMPR11[16] , 
        \R_DATA_TEMPR11[15] , \R_DATA_TEMPR11[14] , 
        \R_DATA_TEMPR11[13] , \R_DATA_TEMPR11[12] , 
        \R_DATA_TEMPR11[11] , \R_DATA_TEMPR11[10] , 
        \R_DATA_TEMPR11[9] , \R_DATA_TEMPR11[8] , \R_DATA_TEMPR11[7] , 
        \R_DATA_TEMPR11[6] , \R_DATA_TEMPR11[5] , \R_DATA_TEMPR11[4] , 
        \R_DATA_TEMPR11[3] , \R_DATA_TEMPR11[2] , \R_DATA_TEMPR11[1] , 
        \R_DATA_TEMPR11[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[11][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[2] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[2] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_3 (.A(\R_DATA_TEMPR8[33] ), .B(\R_DATA_TEMPR9[33] ), .C(
        \R_DATA_TEMPR10[33] ), .D(\R_DATA_TEMPR11[33] ), .Y(OR4_3_Y));
    OR4 OR4_200 (.A(\R_DATA_TEMPR12[52] ), .B(\R_DATA_TEMPR13[52] ), 
        .C(\R_DATA_TEMPR14[52] ), .D(\R_DATA_TEMPR15[52] ), .Y(
        OR4_200_Y));
    OR4 \OR4_R_DATA[34]  (.A(OR4_265_Y), .B(OR4_68_Y), .C(OR4_306_Y), 
        .D(OR4_84_Y), .Y(R_DATA[34]));
    OR4 OR4_242 (.A(\R_DATA_TEMPR12[17] ), .B(\R_DATA_TEMPR13[17] ), 
        .C(\R_DATA_TEMPR14[17] ), .D(\R_DATA_TEMPR15[17] ), .Y(
        OR4_242_Y));
    OR4 OR4_180 (.A(\R_DATA_TEMPR8[18] ), .B(\R_DATA_TEMPR9[18] ), .C(
        \R_DATA_TEMPR10[18] ), .D(\R_DATA_TEMPR11[18] ), .Y(OR4_180_Y));
    OR4 OR4_151 (.A(\R_DATA_TEMPR8[71] ), .B(\R_DATA_TEMPR9[71] ), .C(
        \R_DATA_TEMPR10[71] ), .D(\R_DATA_TEMPR11[71] ), .Y(OR4_151_Y));
    OR4 OR4_86 (.A(\R_DATA_TEMPR0[62] ), .B(\R_DATA_TEMPR1[62] ), .C(
        \R_DATA_TEMPR2[62] ), .D(\R_DATA_TEMPR3[62] ), .Y(OR4_86_Y));
    OR4 \OR4_R_DATA[14]  (.A(OR4_192_Y), .B(OR4_309_Y), .C(OR4_227_Y), 
        .D(OR4_4_Y), .Y(R_DATA[14]));
    OR4 \OR4_R_DATA[33]  (.A(OR4_30_Y), .B(OR4_201_Y), .C(OR4_3_Y), .D(
        OR4_260_Y), .Y(R_DATA[33]));
    OR4 OR4_142 (.A(\R_DATA_TEMPR12[53] ), .B(\R_DATA_TEMPR13[53] ), 
        .C(\R_DATA_TEMPR14[53] ), .D(\R_DATA_TEMPR15[53] ), .Y(
        OR4_142_Y));
    OR4 \OR4_R_DATA[13]  (.A(OR4_277_Y), .B(OR4_113_Y), .C(OR4_248_Y), 
        .D(OR4_181_Y), .Y(R_DATA[13]));
    OR4 \OR4_R_DATA[68]  (.A(OR4_205_Y), .B(OR4_278_Y), .C(OR4_178_Y), 
        .D(OR4_89_Y), .Y(R_DATA[68]));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%7%1%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C1 (.A_DOUT({
        \R_DATA_TEMPR7[79] , \R_DATA_TEMPR7[78] , \R_DATA_TEMPR7[77] , 
        \R_DATA_TEMPR7[76] , \R_DATA_TEMPR7[75] , \R_DATA_TEMPR7[74] , 
        \R_DATA_TEMPR7[73] , \R_DATA_TEMPR7[72] , \R_DATA_TEMPR7[71] , 
        \R_DATA_TEMPR7[70] , \R_DATA_TEMPR7[69] , \R_DATA_TEMPR7[68] , 
        \R_DATA_TEMPR7[67] , \R_DATA_TEMPR7[66] , \R_DATA_TEMPR7[65] , 
        \R_DATA_TEMPR7[64] , \R_DATA_TEMPR7[63] , \R_DATA_TEMPR7[62] , 
        \R_DATA_TEMPR7[61] , \R_DATA_TEMPR7[60] }), .B_DOUT({
        \R_DATA_TEMPR7[59] , \R_DATA_TEMPR7[58] , \R_DATA_TEMPR7[57] , 
        \R_DATA_TEMPR7[56] , \R_DATA_TEMPR7[55] , \R_DATA_TEMPR7[54] , 
        \R_DATA_TEMPR7[53] , \R_DATA_TEMPR7[52] , \R_DATA_TEMPR7[51] , 
        \R_DATA_TEMPR7[50] , \R_DATA_TEMPR7[49] , \R_DATA_TEMPR7[48] , 
        \R_DATA_TEMPR7[47] , \R_DATA_TEMPR7[46] , \R_DATA_TEMPR7[45] , 
        \R_DATA_TEMPR7[44] , \R_DATA_TEMPR7[43] , \R_DATA_TEMPR7[42] , 
        \R_DATA_TEMPR7[41] , \R_DATA_TEMPR7[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[7][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[1] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[66]  (.A(OR4_17_Y), .B(OR4_96_Y), .C(OR4_44_Y), .D(
        OR4_72_Y), .Y(R_DATA[66]));
    OR4 OR4_319 (.A(\R_DATA_TEMPR12[64] ), .B(\R_DATA_TEMPR13[64] ), 
        .C(\R_DATA_TEMPR14[64] ), .D(\R_DATA_TEMPR15[64] ), .Y(
        OR4_319_Y));
    OR4 OR4_111 (.A(\R_DATA_TEMPR12[19] ), .B(\R_DATA_TEMPR13[19] ), 
        .C(\R_DATA_TEMPR14[19] ), .D(\R_DATA_TEMPR15[19] ), .Y(
        OR4_111_Y));
    OR4 \OR4_R_DATA[51]  (.A(OR4_158_Y), .B(OR4_129_Y), .C(OR4_26_Y), 
        .D(OR4_67_Y), .Y(R_DATA[51]));
    OR4 OR4_268 (.A(\R_DATA_TEMPR4[3] ), .B(\R_DATA_TEMPR5[3] ), .C(
        \R_DATA_TEMPR6[3] ), .D(\R_DATA_TEMPR7[3] ), .Y(OR4_268_Y));
    OR4 OR4_226 (.A(\R_DATA_TEMPR0[50] ), .B(\R_DATA_TEMPR1[50] ), .C(
        \R_DATA_TEMPR2[50] ), .D(\R_DATA_TEMPR3[50] ), .Y(OR4_226_Y));
    OR4 OR4_124 (.A(\R_DATA_TEMPR8[22] ), .B(\R_DATA_TEMPR9[22] ), .C(
        \R_DATA_TEMPR10[22] ), .D(\R_DATA_TEMPR11[22] ), .Y(OR4_124_Y));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%10%0%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C0 (.A_DOUT({
        \R_DATA_TEMPR10[39] , \R_DATA_TEMPR10[38] , 
        \R_DATA_TEMPR10[37] , \R_DATA_TEMPR10[36] , 
        \R_DATA_TEMPR10[35] , \R_DATA_TEMPR10[34] , 
        \R_DATA_TEMPR10[33] , \R_DATA_TEMPR10[32] , 
        \R_DATA_TEMPR10[31] , \R_DATA_TEMPR10[30] , 
        \R_DATA_TEMPR10[29] , \R_DATA_TEMPR10[28] , 
        \R_DATA_TEMPR10[27] , \R_DATA_TEMPR10[26] , 
        \R_DATA_TEMPR10[25] , \R_DATA_TEMPR10[24] , 
        \R_DATA_TEMPR10[23] , \R_DATA_TEMPR10[22] , 
        \R_DATA_TEMPR10[21] , \R_DATA_TEMPR10[20] }), .B_DOUT({
        \R_DATA_TEMPR10[19] , \R_DATA_TEMPR10[18] , 
        \R_DATA_TEMPR10[17] , \R_DATA_TEMPR10[16] , 
        \R_DATA_TEMPR10[15] , \R_DATA_TEMPR10[14] , 
        \R_DATA_TEMPR10[13] , \R_DATA_TEMPR10[12] , 
        \R_DATA_TEMPR10[11] , \R_DATA_TEMPR10[10] , 
        \R_DATA_TEMPR10[9] , \R_DATA_TEMPR10[8] , \R_DATA_TEMPR10[7] , 
        \R_DATA_TEMPR10[6] , \R_DATA_TEMPR10[5] , \R_DATA_TEMPR10[4] , 
        \R_DATA_TEMPR10[3] , \R_DATA_TEMPR10[2] , \R_DATA_TEMPR10[1] , 
        \R_DATA_TEMPR10[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[10][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[2] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[2] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[35]  (.A(OR4_136_Y), .B(OR4_125_Y), .C(OR4_272_Y), 
        .D(OR4_244_Y), .Y(R_DATA[35]));
    OR4 OR4_223 (.A(\R_DATA_TEMPR8[64] ), .B(\R_DATA_TEMPR9[64] ), .C(
        \R_DATA_TEMPR10[64] ), .D(\R_DATA_TEMPR11[64] ), .Y(OR4_223_Y));
    OR4 OR4_315 (.A(\R_DATA_TEMPR0[0] ), .B(\R_DATA_TEMPR1[0] ), .C(
        \R_DATA_TEMPR2[0] ), .D(\R_DATA_TEMPR3[0] ), .Y(OR4_315_Y));
    OR4 \OR4_R_DATA[15]  (.A(OR4_62_Y), .B(OR4_43_Y), .C(OR4_199_Y), 
        .D(OR4_160_Y), .Y(R_DATA[15]));
    OR4 \OR4_R_DATA[27]  (.A(OR4_285_Y), .B(OR4_95_Y), .C(OR4_296_Y), 
        .D(OR4_246_Y), .Y(R_DATA[27]));
    OR4 OR4_202 (.A(\R_DATA_TEMPR8[25] ), .B(\R_DATA_TEMPR9[25] ), .C(
        \R_DATA_TEMPR10[25] ), .D(\R_DATA_TEMPR11[25] ), .Y(OR4_202_Y));
    OR4 OR4_276 (.A(\R_DATA_TEMPR0[67] ), .B(\R_DATA_TEMPR1[67] ), .C(
        \R_DATA_TEMPR2[67] ), .D(\R_DATA_TEMPR3[67] ), .Y(OR4_276_Y));
    OR4 OR4_224 (.A(\R_DATA_TEMPR4[0] ), .B(\R_DATA_TEMPR5[0] ), .C(
        \R_DATA_TEMPR6[0] ), .D(\R_DATA_TEMPR7[0] ), .Y(OR4_224_Y));
    OR4 OR4_174 (.A(\R_DATA_TEMPR4[21] ), .B(\R_DATA_TEMPR5[21] ), .C(
        \R_DATA_TEMPR6[21] ), .D(\R_DATA_TEMPR7[21] ), .Y(OR4_174_Y));
    OR4 OR4_291 (.A(\R_DATA_TEMPR8[67] ), .B(\R_DATA_TEMPR9[67] ), .C(
        \R_DATA_TEMPR10[67] ), .D(\R_DATA_TEMPR11[67] ), .Y(OR4_291_Y));
    OR4 OR4_102 (.A(\R_DATA_TEMPR4[39] ), .B(\R_DATA_TEMPR5[39] ), .C(
        \R_DATA_TEMPR6[39] ), .D(\R_DATA_TEMPR7[39] ), .Y(OR4_102_Y));
    OR4 OR4_76 (.A(\R_DATA_TEMPR8[4] ), .B(\R_DATA_TEMPR9[4] ), .C(
        \R_DATA_TEMPR10[4] ), .D(\R_DATA_TEMPR11[4] ), .Y(OR4_76_Y));
    OR4 OR4_273 (.A(\R_DATA_TEMPR8[75] ), .B(\R_DATA_TEMPR9[75] ), .C(
        \R_DATA_TEMPR10[75] ), .D(\R_DATA_TEMPR11[75] ), .Y(OR4_273_Y));
    OR4 OR4_235 (.A(\R_DATA_TEMPR0[53] ), .B(\R_DATA_TEMPR1[53] ), .C(
        \R_DATA_TEMPR2[53] ), .D(\R_DATA_TEMPR3[53] ), .Y(OR4_235_Y));
    OR4 OR4_158 (.A(\R_DATA_TEMPR0[51] ), .B(\R_DATA_TEMPR1[51] ), .C(
        \R_DATA_TEMPR2[51] ), .D(\R_DATA_TEMPR3[51] ), .Y(OR4_158_Y));
    OR4 OR4_23 (.A(\R_DATA_TEMPR0[70] ), .B(\R_DATA_TEMPR1[70] ), .C(
        \R_DATA_TEMPR2[70] ), .D(\R_DATA_TEMPR3[70] ), .Y(OR4_23_Y));
    OR4 OR4_59 (.A(\R_DATA_TEMPR4[32] ), .B(\R_DATA_TEMPR5[32] ), .C(
        \R_DATA_TEMPR6[32] ), .D(\R_DATA_TEMPR7[32] ), .Y(OR4_59_Y));
    OR4 OR4_99 (.A(\R_DATA_TEMPR12[7] ), .B(\R_DATA_TEMPR13[7] ), .C(
        \R_DATA_TEMPR14[7] ), .D(\R_DATA_TEMPR15[7] ), .Y(OR4_99_Y));
    OR4 OR4_186 (.A(\R_DATA_TEMPR12[71] ), .B(\R_DATA_TEMPR13[71] ), 
        .C(\R_DATA_TEMPR14[71] ), .D(\R_DATA_TEMPR15[71] ), .Y(
        OR4_186_Y));
    OR4 OR4_143 (.A(\R_DATA_TEMPR4[8] ), .B(\R_DATA_TEMPR5[8] ), .C(
        \R_DATA_TEMPR6[8] ), .D(\R_DATA_TEMPR7[8] ), .Y(OR4_143_Y));
    OR4 OR4_127 (.A(\R_DATA_TEMPR4[1] ), .B(\R_DATA_TEMPR5[1] ), .C(
        \R_DATA_TEMPR6[1] ), .D(\R_DATA_TEMPR7[1] ), .Y(OR4_127_Y));
    OR4 OR4_274 (.A(\R_DATA_TEMPR0[63] ), .B(\R_DATA_TEMPR1[63] ), .C(
        \R_DATA_TEMPR2[63] ), .D(\R_DATA_TEMPR3[63] ), .Y(OR4_274_Y));
    OR4 OR4_2 (.A(\R_DATA_TEMPR4[55] ), .B(\R_DATA_TEMPR5[55] ), .C(
        \R_DATA_TEMPR6[55] ), .D(\R_DATA_TEMPR7[55] ), .Y(OR4_2_Y));
    OR4 OR4_159 (.A(\R_DATA_TEMPR8[46] ), .B(\R_DATA_TEMPR9[46] ), .C(
        \R_DATA_TEMPR10[46] ), .D(\R_DATA_TEMPR11[46] ), .Y(OR4_159_Y));
    OR4 \OR4_R_DATA[32]  (.A(OR4_164_Y), .B(OR4_59_Y), .C(OR4_206_Y), 
        .D(OR4_311_Y), .Y(R_DATA[32]));
    OR4 OR4_118 (.A(\R_DATA_TEMPR0[8] ), .B(\R_DATA_TEMPR1[8] ), .C(
        \R_DATA_TEMPR2[8] ), .D(\R_DATA_TEMPR3[8] ), .Y(OR4_118_Y));
    OR4 \OR4_R_DATA[12]  (.A(OR4_90_Y), .B(OR4_297_Y), .C(OR4_122_Y), 
        .D(OR4_233_Y), .Y(R_DATA[12]));
    OR4 OR4_38 (.A(\R_DATA_TEMPR4[38] ), .B(\R_DATA_TEMPR5[38] ), .C(
        \R_DATA_TEMPR6[38] ), .D(\R_DATA_TEMPR7[38] ), .Y(OR4_38_Y));
    OR4 OR4_230 (.A(\R_DATA_TEMPR12[62] ), .B(\R_DATA_TEMPR13[62] ), 
        .C(\R_DATA_TEMPR14[62] ), .D(\R_DATA_TEMPR15[62] ), .Y(
        OR4_230_Y));
    OR4 \OR4_R_DATA[20]  (.A(OR4_270_Y), .B(OR4_60_Y), .C(OR4_198_Y), 
        .D(OR4_36_Y), .Y(R_DATA[20]));
    OR4 OR4_155 (.A(\R_DATA_TEMPR0[58] ), .B(\R_DATA_TEMPR1[58] ), .C(
        \R_DATA_TEMPR2[58] ), .D(\R_DATA_TEMPR3[58] ), .Y(OR4_155_Y));
    OR4 OR4_177 (.A(\R_DATA_TEMPR4[76] ), .B(\R_DATA_TEMPR5[76] ), .C(
        \R_DATA_TEMPR6[76] ), .D(\R_DATA_TEMPR7[76] ), .Y(OR4_177_Y));
    OR4 OR4_119 (.A(\R_DATA_TEMPR12[44] ), .B(\R_DATA_TEMPR13[44] ), 
        .C(\R_DATA_TEMPR14[44] ), .D(\R_DATA_TEMPR15[44] ), .Y(
        OR4_119_Y));
    OR4 \OR4_R_DATA[78]  (.A(OR4_281_Y), .B(OR4_39_Y), .C(OR4_261_Y), 
        .D(OR4_172_Y), .Y(R_DATA[78]));
    OR4 \OR4_R_DATA[76]  (.A(OR4_106_Y), .B(OR4_177_Y), .C(OR4_131_Y), 
        .D(OR4_153_Y), .Y(R_DATA[76]));
    OR4 OR4_15 (.A(\R_DATA_TEMPR4[69] ), .B(\R_DATA_TEMPR5[69] ), .C(
        \R_DATA_TEMPR6[69] ), .D(\R_DATA_TEMPR7[69] ), .Y(OR4_15_Y));
    OR4 OR4_65 (.A(\R_DATA_TEMPR0[29] ), .B(\R_DATA_TEMPR1[29] ), .C(
        \R_DATA_TEMPR2[29] ), .D(\R_DATA_TEMPR3[29] ), .Y(OR4_65_Y));
    OR4 \OR4_R_DATA[54]  (.A(OR4_145_Y), .B(OR4_264_Y), .C(OR4_184_Y), 
        .D(OR4_283_Y), .Y(R_DATA[54]));
    OR4 OR4_82 (.A(\R_DATA_TEMPR4[48] ), .B(\R_DATA_TEMPR5[48] ), .C(
        \R_DATA_TEMPR6[48] ), .D(\R_DATA_TEMPR7[48] ), .Y(OR4_82_Y));
    OR4 \OR4_R_DATA[53]  (.A(OR4_235_Y), .B(OR4_75_Y), .C(OR4_213_Y), 
        .D(OR4_142_Y), .Y(R_DATA[53]));
    OR4 OR4_115 (.A(\R_DATA_TEMPR4[23] ), .B(\R_DATA_TEMPR5[23] ), .C(
        \R_DATA_TEMPR6[23] ), .D(\R_DATA_TEMPR7[23] ), .Y(OR4_115_Y));
    OR4 OR4_259 (.A(\R_DATA_TEMPR8[38] ), .B(\R_DATA_TEMPR9[38] ), .C(
        \R_DATA_TEMPR10[38] ), .D(\R_DATA_TEMPR11[38] ), .Y(OR4_259_Y));
    OR4 OR4_160 (.A(\R_DATA_TEMPR12[15] ), .B(\R_DATA_TEMPR13[15] ), 
        .C(\R_DATA_TEMPR14[15] ), .D(\R_DATA_TEMPR15[15] ), .Y(
        OR4_160_Y));
    OR4 OR4_103 (.A(\R_DATA_TEMPR4[79] ), .B(\R_DATA_TEMPR5[79] ), .C(
        \R_DATA_TEMPR6[79] ), .D(\R_DATA_TEMPR7[79] ), .Y(OR4_103_Y));
    OR4 OR4_11 (.A(\R_DATA_TEMPR4[50] ), .B(\R_DATA_TEMPR5[50] ), .C(
        \R_DATA_TEMPR6[50] ), .D(\R_DATA_TEMPR7[50] ), .Y(OR4_11_Y));
    OR4 OR4_61 (.A(\R_DATA_TEMPR4[72] ), .B(\R_DATA_TEMPR5[72] ), .C(
        \R_DATA_TEMPR6[72] ), .D(\R_DATA_TEMPR7[72] ), .Y(OR4_61_Y));
    OR4 OR4_228 (.A(\R_DATA_TEMPR8[24] ), .B(\R_DATA_TEMPR9[24] ), .C(
        \R_DATA_TEMPR10[24] ), .D(\R_DATA_TEMPR11[24] ), .Y(OR4_228_Y));
    OR4 OR4_87 (.A(\R_DATA_TEMPR8[47] ), .B(\R_DATA_TEMPR9[47] ), .C(
        \R_DATA_TEMPR10[47] ), .D(\R_DATA_TEMPR11[47] ), .Y(OR4_87_Y));
    OR4 \OR4_R_DATA[1]  (.A(OR4_247_Y), .B(OR4_127_Y), .C(OR4_150_Y), 
        .D(OR4_1_Y), .Y(R_DATA[1]));
    OR4 OR4_49 (.A(\R_DATA_TEMPR4[60] ), .B(\R_DATA_TEMPR5[60] ), .C(
        \R_DATA_TEMPR6[60] ), .D(\R_DATA_TEMPR7[60] ), .Y(OR4_49_Y));
    OR4 OR4_219 (.A(\R_DATA_TEMPR8[59] ), .B(\R_DATA_TEMPR9[59] ), .C(
        \R_DATA_TEMPR10[59] ), .D(\R_DATA_TEMPR11[59] ), .Y(OR4_219_Y));
    OR4 \OR4_R_DATA[55]  (.A(OR4_13_Y), .B(OR4_2_Y), .C(OR4_148_Y), .D(
        OR4_123_Y), .Y(R_DATA[55]));
    OR4 OR4_303 (.A(\R_DATA_TEMPR4[64] ), .B(\R_DATA_TEMPR5[64] ), .C(
        \R_DATA_TEMPR6[64] ), .D(\R_DATA_TEMPR7[64] ), .Y(OR4_303_Y));
    OR4 OR4_232 (.A(\R_DATA_TEMPR8[42] ), .B(\R_DATA_TEMPR9[42] ), .C(
        \R_DATA_TEMPR10[42] ), .D(\R_DATA_TEMPR11[42] ), .Y(OR4_232_Y));
    OR4 OR4_278 (.A(\R_DATA_TEMPR4[68] ), .B(\R_DATA_TEMPR5[68] ), .C(
        \R_DATA_TEMPR6[68] ), .D(\R_DATA_TEMPR7[68] ), .Y(OR4_278_Y));
    OR4 OR4_132 (.A(\R_DATA_TEMPR4[30] ), .B(\R_DATA_TEMPR5[30] ), .C(
        \R_DATA_TEMPR6[30] ), .D(\R_DATA_TEMPR7[30] ), .Y(OR4_132_Y));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%15%1%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C1 (.A_DOUT({
        \R_DATA_TEMPR15[79] , \R_DATA_TEMPR15[78] , 
        \R_DATA_TEMPR15[77] , \R_DATA_TEMPR15[76] , 
        \R_DATA_TEMPR15[75] , \R_DATA_TEMPR15[74] , 
        \R_DATA_TEMPR15[73] , \R_DATA_TEMPR15[72] , 
        \R_DATA_TEMPR15[71] , \R_DATA_TEMPR15[70] , 
        \R_DATA_TEMPR15[69] , \R_DATA_TEMPR15[68] , 
        \R_DATA_TEMPR15[67] , \R_DATA_TEMPR15[66] , 
        \R_DATA_TEMPR15[65] , \R_DATA_TEMPR15[64] , 
        \R_DATA_TEMPR15[63] , \R_DATA_TEMPR15[62] , 
        \R_DATA_TEMPR15[61] , \R_DATA_TEMPR15[60] }), .B_DOUT({
        \R_DATA_TEMPR15[59] , \R_DATA_TEMPR15[58] , 
        \R_DATA_TEMPR15[57] , \R_DATA_TEMPR15[56] , 
        \R_DATA_TEMPR15[55] , \R_DATA_TEMPR15[54] , 
        \R_DATA_TEMPR15[53] , \R_DATA_TEMPR15[52] , 
        \R_DATA_TEMPR15[51] , \R_DATA_TEMPR15[50] , 
        \R_DATA_TEMPR15[49] , \R_DATA_TEMPR15[48] , 
        \R_DATA_TEMPR15[47] , \R_DATA_TEMPR15[46] , 
        \R_DATA_TEMPR15[45] , \R_DATA_TEMPR15[44] , 
        \R_DATA_TEMPR15[43] , \R_DATA_TEMPR15[42] , 
        \R_DATA_TEMPR15[41] , \R_DATA_TEMPR15[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[15][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[3] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[8]  (.A(OR4_118_Y), .B(OR4_143_Y), .C(OR4_74_Y), 
        .D(OR4_204_Y), .Y(R_DATA[8]));
    OR4 OR4_72 (.A(\R_DATA_TEMPR12[66] ), .B(\R_DATA_TEMPR13[66] ), .C(
        \R_DATA_TEMPR14[66] ), .D(\R_DATA_TEMPR15[66] ), .Y(OR4_72_Y));
    OR4 OR4_241 (.A(\R_DATA_TEMPR4[2] ), .B(\R_DATA_TEMPR5[2] ), .C(
        \R_DATA_TEMPR6[2] ), .D(\R_DATA_TEMPR7[2] ), .Y(OR4_241_Y));
    OR4 OR4_285 (.A(\R_DATA_TEMPR0[27] ), .B(\R_DATA_TEMPR1[27] ), .C(
        \R_DATA_TEMPR2[27] ), .D(\R_DATA_TEMPR3[27] ), .Y(OR4_285_Y));
    OR4 OR4_28 (.A(\R_DATA_TEMPR12[47] ), .B(\R_DATA_TEMPR13[47] ), .C(
        \R_DATA_TEMPR14[47] ), .D(\R_DATA_TEMPR15[47] ), .Y(OR4_28_Y));
    OR4 OR4_54 (.A(\R_DATA_TEMPR8[26] ), .B(\R_DATA_TEMPR9[26] ), .C(
        \R_DATA_TEMPR10[26] ), .D(\R_DATA_TEMPR11[26] ), .Y(OR4_54_Y));
    CFG3 #( .INIT(8'h40) )  \CFG3_BLKX2[1]  (.A(W_ADDR[12]), .B(
        W_ADDR[11]), .C(W_EN), .Y(\BLKX2[1] ));
    OR4 OR4_94 (.A(\R_DATA_TEMPR12[18] ), .B(\R_DATA_TEMPR13[18] ), .C(
        \R_DATA_TEMPR14[18] ), .D(\R_DATA_TEMPR15[18] ), .Y(OR4_94_Y));
    OR4 OR4_77 (.A(\R_DATA_TEMPR0[43] ), .B(\R_DATA_TEMPR1[43] ), .C(
        \R_DATA_TEMPR2[43] ), .D(\R_DATA_TEMPR3[43] ), .Y(OR4_77_Y));
    OR4 \OR4_R_DATA[52]  (.A(OR4_42_Y), .B(OR4_257_Y), .C(OR4_83_Y), 
        .D(OR4_200_Y), .Y(R_DATA[52]));
    OR4 OR4_166 (.A(\R_DATA_TEMPR4[61] ), .B(\R_DATA_TEMPR5[61] ), .C(
        \R_DATA_TEMPR6[61] ), .D(\R_DATA_TEMPR7[61] ), .Y(OR4_166_Y));
    CFG3 #( .INIT(8'h80) )  \CFG3_BLKX2[3]  (.A(W_ADDR[12]), .B(
        W_ADDR[11]), .C(W_EN), .Y(\BLKX2[3] ));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%1%0%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C0 (.A_DOUT({
        \R_DATA_TEMPR1[39] , \R_DATA_TEMPR1[38] , \R_DATA_TEMPR1[37] , 
        \R_DATA_TEMPR1[36] , \R_DATA_TEMPR1[35] , \R_DATA_TEMPR1[34] , 
        \R_DATA_TEMPR1[33] , \R_DATA_TEMPR1[32] , \R_DATA_TEMPR1[31] , 
        \R_DATA_TEMPR1[30] , \R_DATA_TEMPR1[29] , \R_DATA_TEMPR1[28] , 
        \R_DATA_TEMPR1[27] , \R_DATA_TEMPR1[26] , \R_DATA_TEMPR1[25] , 
        \R_DATA_TEMPR1[24] , \R_DATA_TEMPR1[23] , \R_DATA_TEMPR1[22] , 
        \R_DATA_TEMPR1[21] , \R_DATA_TEMPR1[20] }), .B_DOUT({
        \R_DATA_TEMPR1[19] , \R_DATA_TEMPR1[18] , \R_DATA_TEMPR1[17] , 
        \R_DATA_TEMPR1[16] , \R_DATA_TEMPR1[15] , \R_DATA_TEMPR1[14] , 
        \R_DATA_TEMPR1[13] , \R_DATA_TEMPR1[12] , \R_DATA_TEMPR1[11] , 
        \R_DATA_TEMPR1[10] , \R_DATA_TEMPR1[9] , \R_DATA_TEMPR1[8] , 
        \R_DATA_TEMPR1[7] , \R_DATA_TEMPR1[6] , \R_DATA_TEMPR1[5] , 
        \R_DATA_TEMPR1[4] , \R_DATA_TEMPR1[3] , \R_DATA_TEMPR1[2] , 
        \R_DATA_TEMPR1[1] , \R_DATA_TEMPR1[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[1][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[0] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_280 (.A(\R_DATA_TEMPR0[23] ), .B(\R_DATA_TEMPR1[23] ), .C(
        \R_DATA_TEMPR2[23] ), .D(\R_DATA_TEMPR3[23] ), .Y(OR4_280_Y));
    INV \INVBLKX0[0]  (.A(W_ADDR[9]), .Y(\BLKX0[0] ));
    OR4 OR4_36 (.A(\R_DATA_TEMPR12[20] ), .B(\R_DATA_TEMPR13[20] ), .C(
        \R_DATA_TEMPR14[20] ), .D(\R_DATA_TEMPR15[20] ), .Y(OR4_36_Y));
    OR4 OR4_256 (.A(\R_DATA_TEMPR4[5] ), .B(\R_DATA_TEMPR5[5] ), .C(
        \R_DATA_TEMPR6[5] ), .D(\R_DATA_TEMPR7[5] ), .Y(OR4_256_Y));
    OR4 OR4_201 (.A(\R_DATA_TEMPR4[33] ), .B(\R_DATA_TEMPR5[33] ), .C(
        \R_DATA_TEMPR6[33] ), .D(\R_DATA_TEMPR7[33] ), .Y(OR4_201_Y));
    OR4 OR4_154 (.A(\R_DATA_TEMPR12[40] ), .B(\R_DATA_TEMPR13[40] ), 
        .C(\R_DATA_TEMPR14[40] ), .D(\R_DATA_TEMPR15[40] ), .Y(
        OR4_154_Y));
    OR4 OR4_133 (.A(\R_DATA_TEMPR4[70] ), .B(\R_DATA_TEMPR5[70] ), .C(
        \R_DATA_TEMPR6[70] ), .D(\R_DATA_TEMPR7[70] ), .Y(OR4_133_Y));
    OR4 OR4_317 (.A(\R_DATA_TEMPR12[37] ), .B(\R_DATA_TEMPR13[37] ), 
        .C(\R_DATA_TEMPR14[37] ), .D(\R_DATA_TEMPR15[37] ), .Y(
        OR4_317_Y));
    OR4 OR4_253 (.A(\R_DATA_TEMPR8[19] ), .B(\R_DATA_TEMPR9[19] ), .C(
        \R_DATA_TEMPR10[19] ), .D(\R_DATA_TEMPR11[19] ), .Y(OR4_253_Y));
    OR4 \OR4_R_DATA[49]  (.A(OR4_170_Y), .B(OR4_135_Y), .C(OR4_40_Y), 
        .D(OR4_225_Y), .Y(R_DATA[49]));
    OR4 OR4_50 (.A(\R_DATA_TEMPR8[16] ), .B(\R_DATA_TEMPR9[16] ), .C(
        \R_DATA_TEMPR10[16] ), .D(\R_DATA_TEMPR11[16] ), .Y(OR4_50_Y));
    OR4 OR4_120 (.A(\R_DATA_TEMPR12[30] ), .B(\R_DATA_TEMPR13[30] ), 
        .C(\R_DATA_TEMPR14[30] ), .D(\R_DATA_TEMPR15[30] ), .Y(
        OR4_120_Y));
    OR4 OR4_90 (.A(\R_DATA_TEMPR0[12] ), .B(\R_DATA_TEMPR1[12] ), .C(
        \R_DATA_TEMPR2[12] ), .D(\R_DATA_TEMPR3[12] ), .Y(OR4_90_Y));
    OR4 OR4_216 (.A(\R_DATA_TEMPR12[48] ), .B(\R_DATA_TEMPR13[48] ), 
        .C(\R_DATA_TEMPR14[48] ), .D(\R_DATA_TEMPR15[48] ), .Y(
        OR4_216_Y));
    OR4 OR4_114 (.A(\R_DATA_TEMPR0[5] ), .B(\R_DATA_TEMPR1[5] ), .C(
        \R_DATA_TEMPR2[5] ), .D(\R_DATA_TEMPR3[5] ), .Y(OR4_114_Y));
    OR4 OR4_254 (.A(\R_DATA_TEMPR4[71] ), .B(\R_DATA_TEMPR5[71] ), .C(
        \R_DATA_TEMPR6[71] ), .D(\R_DATA_TEMPR7[71] ), .Y(OR4_254_Y));
    OR4 OR4_213 (.A(\R_DATA_TEMPR8[53] ), .B(\R_DATA_TEMPR9[53] ), .C(
        \R_DATA_TEMPR10[53] ), .D(\R_DATA_TEMPR11[53] ), .Y(OR4_213_Y));
    OR4 OR4_44 (.A(\R_DATA_TEMPR8[66] ), .B(\R_DATA_TEMPR9[66] ), .C(
        \R_DATA_TEMPR10[66] ), .D(\R_DATA_TEMPR11[66] ), .Y(OR4_44_Y));
    OR4 OR4_297 (.A(\R_DATA_TEMPR4[12] ), .B(\R_DATA_TEMPR5[12] ), .C(
        \R_DATA_TEMPR6[12] ), .D(\R_DATA_TEMPR7[12] ), .Y(OR4_297_Y));
    OR4 OR4_170 (.A(\R_DATA_TEMPR0[49] ), .B(\R_DATA_TEMPR1[49] ), .C(
        \R_DATA_TEMPR2[49] ), .D(\R_DATA_TEMPR3[49] ), .Y(OR4_170_Y));
    OR4 \OR4_R_DATA[61]  (.A(OR4_209_Y), .B(OR4_166_Y), .C(OR4_70_Y), 
        .D(OR4_104_Y), .Y(R_DATA[61]));
    OR4 \OR4_R_DATA[4]  (.A(OR4_239_Y), .B(OR4_162_Y), .C(OR4_76_Y), 
        .D(OR4_12_Y), .Y(R_DATA[4]));
    CFG3 #( .INIT(8'h20) )  \CFG3_BLKY2[2]  (.A(R_ADDR[12]), .B(
        R_ADDR[11]), .C(R_EN), .Y(\BLKY2[2] ));
    INV \INVBLKX1[0]  (.A(W_ADDR[10]), .Y(\BLKX1[0] ));
    OR4 OR4_282 (.A(\R_DATA_TEMPR0[17] ), .B(\R_DATA_TEMPR1[17] ), .C(
        \R_DATA_TEMPR2[17] ), .D(\R_DATA_TEMPR3[17] ), .Y(OR4_282_Y));
    OR4 OR4_214 (.A(\R_DATA_TEMPR4[47] ), .B(\R_DATA_TEMPR5[47] ), .C(
        \R_DATA_TEMPR6[47] ), .D(\R_DATA_TEMPR7[47] ), .Y(OR4_214_Y));
    OR4 OR4_157 (.A(\R_DATA_TEMPR12[65] ), .B(\R_DATA_TEMPR13[65] ), 
        .C(\R_DATA_TEMPR14[65] ), .D(\R_DATA_TEMPR15[65] ), .Y(
        OR4_157_Y));
    INV \INVBLKY0[0]  (.A(R_ADDR[9]), .Y(\BLKY0[0] ));
    OR4 OR4_182 (.A(\R_DATA_TEMPR8[28] ), .B(\R_DATA_TEMPR9[28] ), .C(
        \R_DATA_TEMPR10[28] ), .D(\R_DATA_TEMPR11[28] ), .Y(OR4_182_Y));
    OR4 OR4_310 (.A(\R_DATA_TEMPR4[24] ), .B(\R_DATA_TEMPR5[24] ), .C(
        \R_DATA_TEMPR6[24] ), .D(\R_DATA_TEMPR7[24] ), .Y(OR4_310_Y));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%2%1%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C1 (.A_DOUT({
        \R_DATA_TEMPR2[79] , \R_DATA_TEMPR2[78] , \R_DATA_TEMPR2[77] , 
        \R_DATA_TEMPR2[76] , \R_DATA_TEMPR2[75] , \R_DATA_TEMPR2[74] , 
        \R_DATA_TEMPR2[73] , \R_DATA_TEMPR2[72] , \R_DATA_TEMPR2[71] , 
        \R_DATA_TEMPR2[70] , \R_DATA_TEMPR2[69] , \R_DATA_TEMPR2[68] , 
        \R_DATA_TEMPR2[67] , \R_DATA_TEMPR2[66] , \R_DATA_TEMPR2[65] , 
        \R_DATA_TEMPR2[64] , \R_DATA_TEMPR2[63] , \R_DATA_TEMPR2[62] , 
        \R_DATA_TEMPR2[61] , \R_DATA_TEMPR2[60] }), .B_DOUT({
        \R_DATA_TEMPR2[59] , \R_DATA_TEMPR2[58] , \R_DATA_TEMPR2[57] , 
        \R_DATA_TEMPR2[56] , \R_DATA_TEMPR2[55] , \R_DATA_TEMPR2[54] , 
        \R_DATA_TEMPR2[53] , \R_DATA_TEMPR2[52] , \R_DATA_TEMPR2[51] , 
        \R_DATA_TEMPR2[50] , \R_DATA_TEMPR2[49] , \R_DATA_TEMPR2[48] , 
        \R_DATA_TEMPR2[47] , \R_DATA_TEMPR2[46] , \R_DATA_TEMPR2[45] , 
        \R_DATA_TEMPR2[44] , \R_DATA_TEMPR2[43] , \R_DATA_TEMPR2[42] , 
        \R_DATA_TEMPR2[41] , \R_DATA_TEMPR2[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[2][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[10], \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[0] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%4%0%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C0 (.A_DOUT({
        \R_DATA_TEMPR4[39] , \R_DATA_TEMPR4[38] , \R_DATA_TEMPR4[37] , 
        \R_DATA_TEMPR4[36] , \R_DATA_TEMPR4[35] , \R_DATA_TEMPR4[34] , 
        \R_DATA_TEMPR4[33] , \R_DATA_TEMPR4[32] , \R_DATA_TEMPR4[31] , 
        \R_DATA_TEMPR4[30] , \R_DATA_TEMPR4[29] , \R_DATA_TEMPR4[28] , 
        \R_DATA_TEMPR4[27] , \R_DATA_TEMPR4[26] , \R_DATA_TEMPR4[25] , 
        \R_DATA_TEMPR4[24] , \R_DATA_TEMPR4[23] , \R_DATA_TEMPR4[22] , 
        \R_DATA_TEMPR4[21] , \R_DATA_TEMPR4[20] }), .B_DOUT({
        \R_DATA_TEMPR4[19] , \R_DATA_TEMPR4[18] , \R_DATA_TEMPR4[17] , 
        \R_DATA_TEMPR4[16] , \R_DATA_TEMPR4[15] , \R_DATA_TEMPR4[14] , 
        \R_DATA_TEMPR4[13] , \R_DATA_TEMPR4[12] , \R_DATA_TEMPR4[11] , 
        \R_DATA_TEMPR4[10] , \R_DATA_TEMPR4[9] , \R_DATA_TEMPR4[8] , 
        \R_DATA_TEMPR4[7] , \R_DATA_TEMPR4[6] , \R_DATA_TEMPR4[5] , 
        \R_DATA_TEMPR4[4] , \R_DATA_TEMPR4[3] , \R_DATA_TEMPR4[2] , 
        \R_DATA_TEMPR4[1] , \R_DATA_TEMPR4[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[4][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[1] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_117 (.A(\R_DATA_TEMPR8[3] ), .B(\R_DATA_TEMPR9[3] ), .C(
        \R_DATA_TEMPR10[3] ), .D(\R_DATA_TEMPR11[3] ), .Y(OR4_117_Y));
    OR4 \OR4_R_DATA[28]  (.A(OR4_212_Y), .B(OR4_290_Y), .C(OR4_182_Y), 
        .D(OR4_97_Y), .Y(R_DATA[28]));
    OR4 OR4_265 (.A(\R_DATA_TEMPR0[34] ), .B(\R_DATA_TEMPR1[34] ), .C(
        \R_DATA_TEMPR2[34] ), .D(\R_DATA_TEMPR3[34] ), .Y(OR4_265_Y));
    OR4 \OR4_R_DATA[26]  (.A(OR4_21_Y), .B(OR4_100_Y), .C(OR4_54_Y), 
        .D(OR4_80_Y), .Y(R_DATA[26]));
    OR4 OR4_26 (.A(\R_DATA_TEMPR8[51] ), .B(\R_DATA_TEMPR9[51] ), .C(
        \R_DATA_TEMPR10[51] ), .D(\R_DATA_TEMPR11[51] ), .Y(OR4_26_Y));
    OR4 OR4_126 (.A(\R_DATA_TEMPR4[75] ), .B(\R_DATA_TEMPR5[75] ), .C(
        \R_DATA_TEMPR6[75] ), .D(\R_DATA_TEMPR7[75] ), .Y(OR4_126_Y));
    OR4 OR4_40 (.A(\R_DATA_TEMPR8[49] ), .B(\R_DATA_TEMPR9[49] ), .C(
        \R_DATA_TEMPR10[49] ), .D(\R_DATA_TEMPR11[49] ), .Y(OR4_40_Y));
    OR4 OR4_85 (.A(\R_DATA_TEMPR12[74] ), .B(\R_DATA_TEMPR13[74] ), .C(
        \R_DATA_TEMPR14[74] ), .D(\R_DATA_TEMPR15[74] ), .Y(OR4_85_Y));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%6%1%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C1 (.A_DOUT({
        \R_DATA_TEMPR6[79] , \R_DATA_TEMPR6[78] , \R_DATA_TEMPR6[77] , 
        \R_DATA_TEMPR6[76] , \R_DATA_TEMPR6[75] , \R_DATA_TEMPR6[74] , 
        \R_DATA_TEMPR6[73] , \R_DATA_TEMPR6[72] , \R_DATA_TEMPR6[71] , 
        \R_DATA_TEMPR6[70] , \R_DATA_TEMPR6[69] , \R_DATA_TEMPR6[68] , 
        \R_DATA_TEMPR6[67] , \R_DATA_TEMPR6[66] , \R_DATA_TEMPR6[65] , 
        \R_DATA_TEMPR6[64] , \R_DATA_TEMPR6[63] , \R_DATA_TEMPR6[62] , 
        \R_DATA_TEMPR6[61] , \R_DATA_TEMPR6[60] }), .B_DOUT({
        \R_DATA_TEMPR6[59] , \R_DATA_TEMPR6[58] , \R_DATA_TEMPR6[57] , 
        \R_DATA_TEMPR6[56] , \R_DATA_TEMPR6[55] , \R_DATA_TEMPR6[54] , 
        \R_DATA_TEMPR6[53] , \R_DATA_TEMPR6[52] , \R_DATA_TEMPR6[51] , 
        \R_DATA_TEMPR6[50] , \R_DATA_TEMPR6[49] , \R_DATA_TEMPR6[48] , 
        \R_DATA_TEMPR6[47] , \R_DATA_TEMPR6[46] , \R_DATA_TEMPR6[45] , 
        \R_DATA_TEMPR6[44] , \R_DATA_TEMPR6[43] , \R_DATA_TEMPR6[42] , 
        \R_DATA_TEMPR6[41] , \R_DATA_TEMPR6[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[6][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[10], \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[1] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_231 (.A(\R_DATA_TEMPR8[2] ), .B(\R_DATA_TEMPR9[2] ), .C(
        \R_DATA_TEMPR10[2] ), .D(\R_DATA_TEMPR11[2] ), .Y(OR4_231_Y));
    OR4 OR4_32 (.A(\R_DATA_TEMPR8[43] ), .B(\R_DATA_TEMPR9[43] ), .C(
        \R_DATA_TEMPR10[43] ), .D(\R_DATA_TEMPR11[43] ), .Y(OR4_32_Y));
    INV \INVBLKY1[0]  (.A(R_ADDR[10]), .Y(\BLKY1[0] ));
    OR4 OR4_81 (.A(\R_DATA_TEMPR0[47] ), .B(\R_DATA_TEMPR1[47] ), .C(
        \R_DATA_TEMPR2[47] ), .D(\R_DATA_TEMPR3[47] ), .Y(OR4_81_Y));
    OR4 OR4_258 (.A(\R_DATA_TEMPR0[7] ), .B(\R_DATA_TEMPR1[7] ), .C(
        \R_DATA_TEMPR2[7] ), .D(\R_DATA_TEMPR3[7] ), .Y(OR4_258_Y));
    OR4 OR4_191 (.A(\R_DATA_TEMPR8[7] ), .B(\R_DATA_TEMPR9[7] ), .C(
        \R_DATA_TEMPR10[7] ), .D(\R_DATA_TEMPR11[7] ), .Y(OR4_191_Y));
    OR4 OR4_176 (.A(\R_DATA_TEMPR4[36] ), .B(\R_DATA_TEMPR5[36] ), .C(
        \R_DATA_TEMPR6[36] ), .D(\R_DATA_TEMPR7[36] ), .Y(OR4_176_Y));
    OR4 OR4_53 (.A(\R_DATA_TEMPR12[2] ), .B(\R_DATA_TEMPR13[2] ), .C(
        \R_DATA_TEMPR14[2] ), .D(\R_DATA_TEMPR15[2] ), .Y(OR4_53_Y));
    OR4 \OR4_R_DATA[47]  (.A(OR4_81_Y), .B(OR4_214_Y), .C(OR4_87_Y), 
        .D(OR4_28_Y), .Y(R_DATA[47]));
    OR4 OR4_93 (.A(\R_DATA_TEMPR4[17] ), .B(\R_DATA_TEMPR5[17] ), .C(
        \R_DATA_TEMPR6[17] ), .D(\R_DATA_TEMPR7[17] ), .Y(OR4_93_Y));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%13%0%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C0 (.A_DOUT({
        \R_DATA_TEMPR13[39] , \R_DATA_TEMPR13[38] , 
        \R_DATA_TEMPR13[37] , \R_DATA_TEMPR13[36] , 
        \R_DATA_TEMPR13[35] , \R_DATA_TEMPR13[34] , 
        \R_DATA_TEMPR13[33] , \R_DATA_TEMPR13[32] , 
        \R_DATA_TEMPR13[31] , \R_DATA_TEMPR13[30] , 
        \R_DATA_TEMPR13[29] , \R_DATA_TEMPR13[28] , 
        \R_DATA_TEMPR13[27] , \R_DATA_TEMPR13[26] , 
        \R_DATA_TEMPR13[25] , \R_DATA_TEMPR13[24] , 
        \R_DATA_TEMPR13[23] , \R_DATA_TEMPR13[22] , 
        \R_DATA_TEMPR13[21] , \R_DATA_TEMPR13[20] }), .B_DOUT({
        \R_DATA_TEMPR13[19] , \R_DATA_TEMPR13[18] , 
        \R_DATA_TEMPR13[17] , \R_DATA_TEMPR13[16] , 
        \R_DATA_TEMPR13[15] , \R_DATA_TEMPR13[14] , 
        \R_DATA_TEMPR13[13] , \R_DATA_TEMPR13[12] , 
        \R_DATA_TEMPR13[11] , \R_DATA_TEMPR13[10] , 
        \R_DATA_TEMPR13[9] , \R_DATA_TEMPR13[8] , \R_DATA_TEMPR13[7] , 
        \R_DATA_TEMPR13[6] , \R_DATA_TEMPR13[5] , \R_DATA_TEMPR13[4] , 
        \R_DATA_TEMPR13[3] , \R_DATA_TEMPR13[2] , \R_DATA_TEMPR13[1] , 
        \R_DATA_TEMPR13[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[13][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[3] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_260 (.A(\R_DATA_TEMPR12[33] ), .B(\R_DATA_TEMPR13[33] ), 
        .C(\R_DATA_TEMPR14[33] ), .D(\R_DATA_TEMPR15[33] ), .Y(
        OR4_260_Y));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%3%1%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C1 (.A_DOUT({
        \R_DATA_TEMPR3[79] , \R_DATA_TEMPR3[78] , \R_DATA_TEMPR3[77] , 
        \R_DATA_TEMPR3[76] , \R_DATA_TEMPR3[75] , \R_DATA_TEMPR3[74] , 
        \R_DATA_TEMPR3[73] , \R_DATA_TEMPR3[72] , \R_DATA_TEMPR3[71] , 
        \R_DATA_TEMPR3[70] , \R_DATA_TEMPR3[69] , \R_DATA_TEMPR3[68] , 
        \R_DATA_TEMPR3[67] , \R_DATA_TEMPR3[66] , \R_DATA_TEMPR3[65] , 
        \R_DATA_TEMPR3[64] , \R_DATA_TEMPR3[63] , \R_DATA_TEMPR3[62] , 
        \R_DATA_TEMPR3[61] , \R_DATA_TEMPR3[60] }), .B_DOUT({
        \R_DATA_TEMPR3[59] , \R_DATA_TEMPR3[58] , \R_DATA_TEMPR3[57] , 
        \R_DATA_TEMPR3[56] , \R_DATA_TEMPR3[55] , \R_DATA_TEMPR3[54] , 
        \R_DATA_TEMPR3[53] , \R_DATA_TEMPR3[52] , \R_DATA_TEMPR3[51] , 
        \R_DATA_TEMPR3[50] , \R_DATA_TEMPR3[49] , \R_DATA_TEMPR3[48] , 
        \R_DATA_TEMPR3[47] , \R_DATA_TEMPR3[46] , \R_DATA_TEMPR3[45] , 
        \R_DATA_TEMPR3[44] , \R_DATA_TEMPR3[43] , \R_DATA_TEMPR3[42] , 
        \R_DATA_TEMPR3[41] , \R_DATA_TEMPR3[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[3][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[0] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_183 (.A(\R_DATA_TEMPR12[23] ), .B(\R_DATA_TEMPR13[23] ), 
        .C(\R_DATA_TEMPR14[23] ), .D(\R_DATA_TEMPR15[23] ), .Y(
        OR4_183_Y));
    OR4 \OR4_R_DATA[64]  (.A(OR4_187_Y), .B(OR4_303_Y), .C(OR4_223_Y), 
        .D(OR4_319_Y), .Y(R_DATA[64]));
    OR4 \OR4_R_DATA[71]  (.A(OR4_286_Y), .B(OR4_254_Y), .C(OR4_151_Y), 
        .D(OR4_186_Y), .Y(R_DATA[71]));
    OR4 OR4_218 (.A(\R_DATA_TEMPR12[9] ), .B(\R_DATA_TEMPR13[9] ), .C(
        \R_DATA_TEMPR14[9] ), .D(\R_DATA_TEMPR15[9] ), .Y(OR4_218_Y));
    OR4 OR4_37 (.A(\R_DATA_TEMPR4[65] ), .B(\R_DATA_TEMPR5[65] ), .C(
        \R_DATA_TEMPR6[65] ), .D(\R_DATA_TEMPR7[65] ), .Y(OR4_37_Y));
    OR4 OR4_5 (.A(\R_DATA_TEMPR8[73] ), .B(\R_DATA_TEMPR9[73] ), .C(
        \R_DATA_TEMPR10[73] ), .D(\R_DATA_TEMPR11[73] ), .Y(OR4_5_Y));
    OR4 OR4_9 (.A(\R_DATA_TEMPR8[79] ), .B(\R_DATA_TEMPR9[79] ), .C(
        \R_DATA_TEMPR10[79] ), .D(\R_DATA_TEMPR11[79] ), .Y(OR4_9_Y));
    OR4 \OR4_R_DATA[63]  (.A(OR4_274_Y), .B(OR4_110_Y), .C(OR4_243_Y), 
        .D(OR4_179_Y), .Y(R_DATA[63]));
    OR4 OR4_75 (.A(\R_DATA_TEMPR4[53] ), .B(\R_DATA_TEMPR5[53] ), .C(
        \R_DATA_TEMPR6[53] ), .D(\R_DATA_TEMPR7[53] ), .Y(OR4_75_Y));
    OR4 OR4_304 (.A(\R_DATA_TEMPR8[40] ), .B(\R_DATA_TEMPR9[40] ), .C(
        \R_DATA_TEMPR10[40] ), .D(\R_DATA_TEMPR11[40] ), .Y(OR4_304_Y));
    OR4 OR4_247 (.A(\R_DATA_TEMPR0[1] ), .B(\R_DATA_TEMPR1[1] ), .C(
        \R_DATA_TEMPR2[1] ), .D(\R_DATA_TEMPR3[1] ), .Y(OR4_247_Y));
    OR4 \OR4_R_DATA[65]  (.A(OR4_55_Y), .B(OR4_37_Y), .C(OR4_193_Y), 
        .D(OR4_157_Y), .Y(R_DATA[65]));
    OR4 OR4_71 (.A(\R_DATA_TEMPR12[59] ), .B(\R_DATA_TEMPR13[59] ), .C(
        \R_DATA_TEMPR14[59] ), .D(\R_DATA_TEMPR15[59] ), .Y(OR4_71_Y));
    OR4 OR4_316 (.A(\R_DATA_TEMPR12[50] ), .B(\R_DATA_TEMPR13[50] ), 
        .C(\R_DATA_TEMPR14[50] ), .D(\R_DATA_TEMPR15[50] ), .Y(
        OR4_316_Y));
    OR4 OR4_198 (.A(\R_DATA_TEMPR8[20] ), .B(\R_DATA_TEMPR9[20] ), .C(
        \R_DATA_TEMPR10[20] ), .D(\R_DATA_TEMPR11[20] ), .Y(OR4_198_Y));
    OR4 OR4_262 (.A(\R_DATA_TEMPR12[73] ), .B(\R_DATA_TEMPR13[73] ), 
        .C(\R_DATA_TEMPR14[73] ), .D(\R_DATA_TEMPR15[73] ), .Y(
        OR4_262_Y));
    OR4 OR4_318 (.A(\R_DATA_TEMPR12[77] ), .B(\R_DATA_TEMPR13[77] ), 
        .C(\R_DATA_TEMPR14[77] ), .D(\R_DATA_TEMPR15[77] ), .Y(
        OR4_318_Y));
    OR4 \OR4_R_DATA[40]  (.A(OR4_66_Y), .B(OR4_163_Y), .C(OR4_304_Y), 
        .D(OR4_154_Y), .Y(R_DATA[40]));
    OR4 OR4_301 (.A(\R_DATA_TEMPR0[44] ), .B(\R_DATA_TEMPR1[44] ), .C(
        \R_DATA_TEMPR2[44] ), .D(\R_DATA_TEMPR3[44] ), .Y(OR4_301_Y));
    OR4 OR4_162 (.A(\R_DATA_TEMPR4[4] ), .B(\R_DATA_TEMPR5[4] ), .C(
        \R_DATA_TEMPR6[4] ), .D(\R_DATA_TEMPR7[4] ), .Y(OR4_162_Y));
    OR4 OR4_43 (.A(\R_DATA_TEMPR4[15] ), .B(\R_DATA_TEMPR5[15] ), .C(
        \R_DATA_TEMPR6[15] ), .D(\R_DATA_TEMPR7[15] ), .Y(OR4_43_Y));
    OR4 OR4_225 (.A(\R_DATA_TEMPR12[49] ), .B(\R_DATA_TEMPR13[49] ), 
        .C(\R_DATA_TEMPR14[49] ), .D(\R_DATA_TEMPR15[49] ), .Y(
        OR4_225_Y));
    OR4 OR4_199 (.A(\R_DATA_TEMPR8[15] ), .B(\R_DATA_TEMPR9[15] ), .C(
        \R_DATA_TEMPR10[15] ), .D(\R_DATA_TEMPR11[15] ), .Y(OR4_199_Y));
    OR4 OR4_22 (.A(\R_DATA_TEMPR0[30] ), .B(\R_DATA_TEMPR1[30] ), .C(
        \R_DATA_TEMPR2[30] ), .D(\R_DATA_TEMPR3[30] ), .Y(OR4_22_Y));
    CFG3 #( .INIT(8'h10) )  \CFG3_BLKY2[0]  (.A(R_ADDR[12]), .B(
        R_ADDR[11]), .C(R_EN), .Y(\BLKY2[0] ));
    OR4 OR4_207 (.A(\R_DATA_TEMPR8[72] ), .B(\R_DATA_TEMPR9[72] ), .C(
        \R_DATA_TEMPR10[72] ), .D(\R_DATA_TEMPR11[72] ), .Y(OR4_207_Y));
    OR4 OR4_4 (.A(\R_DATA_TEMPR12[14] ), .B(\R_DATA_TEMPR13[14] ), .C(
        \R_DATA_TEMPR14[14] ), .D(\R_DATA_TEMPR15[14] ), .Y(OR4_4_Y));
    OR4 OR4_195 (.A(\R_DATA_TEMPR12[39] ), .B(\R_DATA_TEMPR13[39] ), 
        .C(\R_DATA_TEMPR14[39] ), .D(\R_DATA_TEMPR15[39] ), .Y(
        OR4_195_Y));
    OR4 OR4_150 (.A(\R_DATA_TEMPR8[1] ), .B(\R_DATA_TEMPR9[1] ), .C(
        \R_DATA_TEMPR10[1] ), .D(\R_DATA_TEMPR11[1] ), .Y(OR4_150_Y));
    OR4 \OR4_R_DATA[62]  (.A(OR4_86_Y), .B(OR4_293_Y), .C(OR4_116_Y), 
        .D(OR4_230_Y), .Y(R_DATA[62]));
    OR4 OR4_275 (.A(\R_DATA_TEMPR12[45] ), .B(\R_DATA_TEMPR13[45] ), 
        .C(\R_DATA_TEMPR14[45] ), .D(\R_DATA_TEMPR15[45] ), .Y(
        OR4_275_Y));
    OR4 OR4_69 (.A(\R_DATA_TEMPR4[74] ), .B(\R_DATA_TEMPR5[74] ), .C(
        \R_DATA_TEMPR6[74] ), .D(\R_DATA_TEMPR7[74] ), .Y(OR4_69_Y));
    OR4 OR4_19 (.A(\R_DATA_TEMPR4[29] ), .B(\R_DATA_TEMPR5[29] ), .C(
        \R_DATA_TEMPR6[29] ), .D(\R_DATA_TEMPR7[29] ), .Y(OR4_19_Y));
    OR4 OR4_27 (.A(\R_DATA_TEMPR12[56] ), .B(\R_DATA_TEMPR13[56] ), .C(
        \R_DATA_TEMPR14[56] ), .D(\R_DATA_TEMPR15[56] ), .Y(OR4_27_Y));
    OR4 \OR4_R_DATA[39]  (.A(OR4_138_Y), .B(OR4_102_Y), .C(OR4_8_Y), 
        .D(OR4_195_Y), .Y(R_DATA[39]));
    OR4 \OR4_R_DATA[74]  (.A(OR4_266_Y), .B(OR4_69_Y), .C(OR4_307_Y), 
        .D(OR4_85_Y), .Y(R_DATA[74]));
    OR4 OR4_281 (.A(\R_DATA_TEMPR0[78] ), .B(\R_DATA_TEMPR1[78] ), .C(
        \R_DATA_TEMPR2[78] ), .D(\R_DATA_TEMPR3[78] ), .Y(OR4_281_Y));
    OR4 \OR4_R_DATA[0]  (.A(OR4_315_Y), .B(OR4_224_Y), .C(OR4_144_Y), 
        .D(OR4_298_Y), .Y(R_DATA[0]));
    OR4 OR4_141 (.A(\R_DATA_TEMPR8[58] ), .B(\R_DATA_TEMPR9[58] ), .C(
        \R_DATA_TEMPR10[58] ), .D(\R_DATA_TEMPR11[58] ), .Y(OR4_141_Y));
    OR4 \OR4_R_DATA[73]  (.A(OR4_31_Y), .B(OR4_203_Y), .C(OR4_5_Y), .D(
        OR4_262_Y), .Y(R_DATA[73]));
    OR4 OR4_220 (.A(\R_DATA_TEMPR4[46] ), .B(\R_DATA_TEMPR5[46] ), .C(
        \R_DATA_TEMPR6[46] ), .D(\R_DATA_TEMPR7[46] ), .Y(OR4_220_Y));
    OR4 \OR4_R_DATA[19]  (.A(OR4_63_Y), .B(OR4_18_Y), .C(OR4_253_Y), 
        .D(OR4_111_Y), .Y(R_DATA[19]));
    OR4 OR4_110 (.A(\R_DATA_TEMPR4[63] ), .B(\R_DATA_TEMPR5[63] ), .C(
        \R_DATA_TEMPR6[63] ), .D(\R_DATA_TEMPR7[63] ), .Y(OR4_110_Y));
    OR4 OR4_58 (.A(\R_DATA_TEMPR4[56] ), .B(\R_DATA_TEMPR5[56] ), .C(
        \R_DATA_TEMPR6[56] ), .D(\R_DATA_TEMPR7[56] ), .Y(OR4_58_Y));
    OR4 OR4_299 (.A(\R_DATA_TEMPR4[22] ), .B(\R_DATA_TEMPR5[22] ), .C(
        \R_DATA_TEMPR6[22] ), .D(\R_DATA_TEMPR7[22] ), .Y(OR4_299_Y));
    OR4 OR4_98 (.A(\R_DATA_TEMPR4[16] ), .B(\R_DATA_TEMPR5[16] ), .C(
        \R_DATA_TEMPR6[16] ), .D(\R_DATA_TEMPR7[16] ), .Y(OR4_98_Y));
    OR4 OR4_163 (.A(\R_DATA_TEMPR4[40] ), .B(\R_DATA_TEMPR5[40] ), .C(
        \R_DATA_TEMPR6[40] ), .D(\R_DATA_TEMPR7[40] ), .Y(OR4_163_Y));
    OR4 OR4_270 (.A(\R_DATA_TEMPR0[20] ), .B(\R_DATA_TEMPR1[20] ), .C(
        \R_DATA_TEMPR2[20] ), .D(\R_DATA_TEMPR3[20] ), .Y(OR4_270_Y));
    OR4 \OR4_R_DATA[75]  (.A(OR4_137_Y), .B(OR4_126_Y), .C(OR4_273_Y), 
        .D(OR4_245_Y), .Y(R_DATA[75]));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%7%0%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C0 (.A_DOUT({
        \R_DATA_TEMPR7[39] , \R_DATA_TEMPR7[38] , \R_DATA_TEMPR7[37] , 
        \R_DATA_TEMPR7[36] , \R_DATA_TEMPR7[35] , \R_DATA_TEMPR7[34] , 
        \R_DATA_TEMPR7[33] , \R_DATA_TEMPR7[32] , \R_DATA_TEMPR7[31] , 
        \R_DATA_TEMPR7[30] , \R_DATA_TEMPR7[29] , \R_DATA_TEMPR7[28] , 
        \R_DATA_TEMPR7[27] , \R_DATA_TEMPR7[26] , \R_DATA_TEMPR7[25] , 
        \R_DATA_TEMPR7[24] , \R_DATA_TEMPR7[23] , \R_DATA_TEMPR7[22] , 
        \R_DATA_TEMPR7[21] , \R_DATA_TEMPR7[20] }), .B_DOUT({
        \R_DATA_TEMPR7[19] , \R_DATA_TEMPR7[18] , \R_DATA_TEMPR7[17] , 
        \R_DATA_TEMPR7[16] , \R_DATA_TEMPR7[15] , \R_DATA_TEMPR7[14] , 
        \R_DATA_TEMPR7[13] , \R_DATA_TEMPR7[12] , \R_DATA_TEMPR7[11] , 
        \R_DATA_TEMPR7[10] , \R_DATA_TEMPR7[9] , \R_DATA_TEMPR7[8] , 
        \R_DATA_TEMPR7[7] , \R_DATA_TEMPR7[6] , \R_DATA_TEMPR7[5] , 
        \R_DATA_TEMPR7[4] , \R_DATA_TEMPR7[3] , \R_DATA_TEMPR7[2] , 
        \R_DATA_TEMPR7[1] , \R_DATA_TEMPR7[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[7][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[1] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_309 (.A(\R_DATA_TEMPR4[14] ), .B(\R_DATA_TEMPR5[14] ), .C(
        \R_DATA_TEMPR6[14] ), .D(\R_DATA_TEMPR7[14] ), .Y(OR4_309_Y));
    OR4 OR4_101 (.A(\R_DATA_TEMPR4[44] ), .B(\R_DATA_TEMPR5[44] ), .C(
        \R_DATA_TEMPR6[44] ), .D(\R_DATA_TEMPR7[44] ), .Y(OR4_101_Y));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%14%1%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C1 (.A_DOUT({
        \R_DATA_TEMPR14[79] , \R_DATA_TEMPR14[78] , 
        \R_DATA_TEMPR14[77] , \R_DATA_TEMPR14[76] , 
        \R_DATA_TEMPR14[75] , \R_DATA_TEMPR14[74] , 
        \R_DATA_TEMPR14[73] , \R_DATA_TEMPR14[72] , 
        \R_DATA_TEMPR14[71] , \R_DATA_TEMPR14[70] , 
        \R_DATA_TEMPR14[69] , \R_DATA_TEMPR14[68] , 
        \R_DATA_TEMPR14[67] , \R_DATA_TEMPR14[66] , 
        \R_DATA_TEMPR14[65] , \R_DATA_TEMPR14[64] , 
        \R_DATA_TEMPR14[63] , \R_DATA_TEMPR14[62] , 
        \R_DATA_TEMPR14[61] , \R_DATA_TEMPR14[60] }), .B_DOUT({
        \R_DATA_TEMPR14[59] , \R_DATA_TEMPR14[58] , 
        \R_DATA_TEMPR14[57] , \R_DATA_TEMPR14[56] , 
        \R_DATA_TEMPR14[55] , \R_DATA_TEMPR14[54] , 
        \R_DATA_TEMPR14[53] , \R_DATA_TEMPR14[52] , 
        \R_DATA_TEMPR14[51] , \R_DATA_TEMPR14[50] , 
        \R_DATA_TEMPR14[49] , \R_DATA_TEMPR14[48] , 
        \R_DATA_TEMPR14[47] , \R_DATA_TEMPR14[46] , 
        \R_DATA_TEMPR14[45] , \R_DATA_TEMPR14[44] , 
        \R_DATA_TEMPR14[43] , \R_DATA_TEMPR14[42] , 
        \R_DATA_TEMPR14[41] , \R_DATA_TEMPR14[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[14][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[10], \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[3] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_222 (.A(\R_DATA_TEMPR12[41] ), .B(\R_DATA_TEMPR13[41] ), 
        .C(\R_DATA_TEMPR14[41] ), .D(\R_DATA_TEMPR15[41] ), .Y(
        OR4_222_Y));
    OR4 OR4_156 (.A(\R_DATA_TEMPR4[45] ), .B(\R_DATA_TEMPR5[45] ), .C(
        \R_DATA_TEMPR6[45] ), .D(\R_DATA_TEMPR7[45] ), .Y(OR4_156_Y));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%2%0%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C0 (.A_DOUT({
        \R_DATA_TEMPR2[39] , \R_DATA_TEMPR2[38] , \R_DATA_TEMPR2[37] , 
        \R_DATA_TEMPR2[36] , \R_DATA_TEMPR2[35] , \R_DATA_TEMPR2[34] , 
        \R_DATA_TEMPR2[33] , \R_DATA_TEMPR2[32] , \R_DATA_TEMPR2[31] , 
        \R_DATA_TEMPR2[30] , \R_DATA_TEMPR2[29] , \R_DATA_TEMPR2[28] , 
        \R_DATA_TEMPR2[27] , \R_DATA_TEMPR2[26] , \R_DATA_TEMPR2[25] , 
        \R_DATA_TEMPR2[24] , \R_DATA_TEMPR2[23] , \R_DATA_TEMPR2[22] , 
        \R_DATA_TEMPR2[21] , \R_DATA_TEMPR2[20] }), .B_DOUT({
        \R_DATA_TEMPR2[19] , \R_DATA_TEMPR2[18] , \R_DATA_TEMPR2[17] , 
        \R_DATA_TEMPR2[16] , \R_DATA_TEMPR2[15] , \R_DATA_TEMPR2[14] , 
        \R_DATA_TEMPR2[13] , \R_DATA_TEMPR2[12] , \R_DATA_TEMPR2[11] , 
        \R_DATA_TEMPR2[10] , \R_DATA_TEMPR2[9] , \R_DATA_TEMPR2[8] , 
        \R_DATA_TEMPR2[7] , \R_DATA_TEMPR2[6] , \R_DATA_TEMPR2[5] , 
        \R_DATA_TEMPR2[4] , \R_DATA_TEMPR2[3] , \R_DATA_TEMPR2[2] , 
        \R_DATA_TEMPR2[1] , \R_DATA_TEMPR2[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[2][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[10], \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[0] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_148 (.A(\R_DATA_TEMPR8[55] ), .B(\R_DATA_TEMPR9[55] ), .C(
        \R_DATA_TEMPR10[55] ), .D(\R_DATA_TEMPR11[55] ), .Y(OR4_148_Y));
    OR4 OR4_305 (.A(\R_DATA_TEMPR4[9] ), .B(\R_DATA_TEMPR5[9] ), .C(
        \R_DATA_TEMPR6[9] ), .D(\R_DATA_TEMPR7[9] ), .Y(OR4_305_Y));
    OR4 OR4_122 (.A(\R_DATA_TEMPR8[12] ), .B(\R_DATA_TEMPR9[12] ), .C(
        \R_DATA_TEMPR10[12] ), .D(\R_DATA_TEMPR11[12] ), .Y(OR4_122_Y));
    OR4 \OR4_R_DATA[2]  (.A(OR4_25_Y), .B(OR4_241_Y), .C(OR4_231_Y), 
        .D(OR4_53_Y), .Y(R_DATA[2]));
    OR4 OR4_116 (.A(\R_DATA_TEMPR8[62] ), .B(\R_DATA_TEMPR9[62] ), .C(
        \R_DATA_TEMPR10[62] ), .D(\R_DATA_TEMPR11[62] ), .Y(OR4_116_Y));
    OR4 OR4_35 (.A(\R_DATA_TEMPR0[77] ), .B(\R_DATA_TEMPR1[77] ), .C(
        \R_DATA_TEMPR2[77] ), .D(\R_DATA_TEMPR3[77] ), .Y(OR4_35_Y));
    OR4 OR4_237 (.A(\R_DATA_TEMPR12[67] ), .B(\R_DATA_TEMPR13[67] ), 
        .C(\R_DATA_TEMPR14[67] ), .D(\R_DATA_TEMPR15[67] ), .Y(
        OR4_237_Y));
    OR4 OR4_149 (.A(\R_DATA_TEMPR8[31] ), .B(\R_DATA_TEMPR9[31] ), .C(
        \R_DATA_TEMPR10[31] ), .D(\R_DATA_TEMPR11[31] ), .Y(OR4_149_Y));
    OR4 \OR4_R_DATA[72]  (.A(OR4_165_Y), .B(OR4_61_Y), .C(OR4_207_Y), 
        .D(OR4_312_Y), .Y(R_DATA[72]));
    OR4 OR4_48 (.A(\R_DATA_TEMPR12[58] ), .B(\R_DATA_TEMPR13[58] ), .C(
        \R_DATA_TEMPR14[58] ), .D(\R_DATA_TEMPR15[58] ), .Y(OR4_48_Y));
    OR4 OR4_272 (.A(\R_DATA_TEMPR8[35] ), .B(\R_DATA_TEMPR9[35] ), .C(
        \R_DATA_TEMPR10[35] ), .D(\R_DATA_TEMPR11[35] ), .Y(OR4_272_Y));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%13%1%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C1 (.A_DOUT({
        \R_DATA_TEMPR13[79] , \R_DATA_TEMPR13[78] , 
        \R_DATA_TEMPR13[77] , \R_DATA_TEMPR13[76] , 
        \R_DATA_TEMPR13[75] , \R_DATA_TEMPR13[74] , 
        \R_DATA_TEMPR13[73] , \R_DATA_TEMPR13[72] , 
        \R_DATA_TEMPR13[71] , \R_DATA_TEMPR13[70] , 
        \R_DATA_TEMPR13[69] , \R_DATA_TEMPR13[68] , 
        \R_DATA_TEMPR13[67] , \R_DATA_TEMPR13[66] , 
        \R_DATA_TEMPR13[65] , \R_DATA_TEMPR13[64] , 
        \R_DATA_TEMPR13[63] , \R_DATA_TEMPR13[62] , 
        \R_DATA_TEMPR13[61] , \R_DATA_TEMPR13[60] }), .B_DOUT({
        \R_DATA_TEMPR13[59] , \R_DATA_TEMPR13[58] , 
        \R_DATA_TEMPR13[57] , \R_DATA_TEMPR13[56] , 
        \R_DATA_TEMPR13[55] , \R_DATA_TEMPR13[54] , 
        \R_DATA_TEMPR13[53] , \R_DATA_TEMPR13[52] , 
        \R_DATA_TEMPR13[51] , \R_DATA_TEMPR13[50] , 
        \R_DATA_TEMPR13[49] , \R_DATA_TEMPR13[48] , 
        \R_DATA_TEMPR13[47] , \R_DATA_TEMPR13[46] , 
        \R_DATA_TEMPR13[45] , \R_DATA_TEMPR13[44] , 
        \R_DATA_TEMPR13[43] , \R_DATA_TEMPR13[42] , 
        \R_DATA_TEMPR13[41] , \R_DATA_TEMPR13[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[13][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[3] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM%8192-8192%80-80%POWER%8%0%TWO-PORT%ECC_EN-0")
         )  LSRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C0 (.A_DOUT({
        \R_DATA_TEMPR8[39] , \R_DATA_TEMPR8[38] , \R_DATA_TEMPR8[37] , 
        \R_DATA_TEMPR8[36] , \R_DATA_TEMPR8[35] , \R_DATA_TEMPR8[34] , 
        \R_DATA_TEMPR8[33] , \R_DATA_TEMPR8[32] , \R_DATA_TEMPR8[31] , 
        \R_DATA_TEMPR8[30] , \R_DATA_TEMPR8[29] , \R_DATA_TEMPR8[28] , 
        \R_DATA_TEMPR8[27] , \R_DATA_TEMPR8[26] , \R_DATA_TEMPR8[25] , 
        \R_DATA_TEMPR8[24] , \R_DATA_TEMPR8[23] , \R_DATA_TEMPR8[22] , 
        \R_DATA_TEMPR8[21] , \R_DATA_TEMPR8[20] }), .B_DOUT({
        \R_DATA_TEMPR8[19] , \R_DATA_TEMPR8[18] , \R_DATA_TEMPR8[17] , 
        \R_DATA_TEMPR8[16] , \R_DATA_TEMPR8[15] , \R_DATA_TEMPR8[14] , 
        \R_DATA_TEMPR8[13] , \R_DATA_TEMPR8[12] , \R_DATA_TEMPR8[11] , 
        \R_DATA_TEMPR8[10] , \R_DATA_TEMPR8[9] , \R_DATA_TEMPR8[8] , 
        \R_DATA_TEMPR8[7] , \R_DATA_TEMPR8[6] , \R_DATA_TEMPR8[5] , 
        \R_DATA_TEMPR8[4] , \R_DATA_TEMPR8[3] , \R_DATA_TEMPR8[2] , 
        \R_DATA_TEMPR8[1] , \R_DATA_TEMPR8[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[8][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[2] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    GND GND_power_inst1 (.Y(GND_power_net1));
    VCC VCC_power_inst1 (.Y(VCC_power_net1));
    
endmodule
